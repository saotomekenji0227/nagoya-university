/*******************/
/* rom8x1024_sim.v */
/*******************/

//                  +----+
//  rom_addr[11:0]->|    |->rom_data[31:0]
//                  +----+

//
// ROM�ε��ҡ��������ߥ�졼������ѡ�
//

module rom8x1024_sim (rom_addr, rom_data);

  input   [11:0]  rom_addr;  // 12-bit ���ɥ쥹���ϥݡ���
  output  [31:0]  rom_data;  // 32-bit �ǡ������ϥݡ���

  reg     [31:0]  data;

  // Wire
  wire     [9:0]  word_addr; // 10-bit address, word

  assign word_addr = rom_addr[9:2];
   
  always @(word_addr) begin
    case (word_addr)
      10'h000: data = 32'he000001c; // 00400000: other type! opcode=56(10)
      10'h001: data = 32'h00000000; // 00400004: SLL, REG[0]<=REG[0]<<0;
      10'h002: data = 32'h00000000; // 00400008: SLL, REG[0]<=REG[0]<<0;
      10'h003: data = 32'h00000000; // 0040000c: SLL, REG[0]<=REG[0]<<0;
      10'h004: data = 32'h00000000; // 00400010: SLL, REG[0]<=REG[0]<<0;
      10'h005: data = 32'h004083d0; // 00400014: R type, unknown. func=16(10)
      10'h006: data = 32'h00000000; // 00400018: SLL, REG[0]<=REG[0]<<0;
      10'h007: data = 32'h00000000; // 0040001c: SLL, REG[0]<=REG[0]<<0;
      10'h008: data = 32'h27bdfee8; // 00400020: ADDIU, REG[29]<=REG[29]+65256(=0x0000fee8);
      10'h009: data = 32'hafbf0114; // 00400024: SW, RAM[REG[29]+276]<=REG[31];
      10'h00a: data = 32'hafbe0110; // 00400028: SW, RAM[REG[29]+272]<=REG[30];
      10'h00b: data = 32'h03a0f021; // 0040002c: ADDU, REG[30]<=REG[29]+REG[0];
      10'h00c: data = 32'h24020048; // 00400030: ADDIU, REG[2]<=REG[0]+72(=0x00000048);
      10'h00d: data = 32'hafc20010; // 00400034: SW, RAM[REG[30]+16]<=REG[2];
      10'h00e: data = 32'h24020045; // 00400038: ADDIU, REG[2]<=REG[0]+69(=0x00000045);
      10'h00f: data = 32'hafc20014; // 0040003c: SW, RAM[REG[30]+20]<=REG[2];
      10'h010: data = 32'h2402004c; // 00400040: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h011: data = 32'hafc20018; // 00400044: SW, RAM[REG[30]+24]<=REG[2];
      10'h012: data = 32'h2402004c; // 00400048: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h013: data = 32'hafc2001c; // 0040004c: SW, RAM[REG[30]+28]<=REG[2];
      10'h014: data = 32'h2402004f; // 00400050: ADDIU, REG[2]<=REG[0]+79(=0x0000004f);
      10'h015: data = 32'hafc20020; // 00400054: SW, RAM[REG[30]+32]<=REG[2];
      10'h016: data = 32'h24020021; // 00400058: ADDIU, REG[2]<=REG[0]+33(=0x00000021);
      10'h017: data = 32'hafc20024; // 0040005c: SW, RAM[REG[30]+36]<=REG[2];
      10'h018: data = 32'h24020021; // 00400060: ADDIU, REG[2]<=REG[0]+33(=0x00000021);
      10'h019: data = 32'hafc20028; // 00400064: SW, RAM[REG[30]+40]<=REG[2];
      10'h01a: data = 32'hafc0002c; // 00400068: SW, RAM[REG[30]+44]<=REG[0];
      10'h01b: data = 32'h27c20010; // 0040006c: ADDIU, REG[2]<=REG[30]+16(=0x00000010);
      10'h01c: data = 32'h00402021; // 00400070: ADDU, REG[4]<=REG[2]+REG[0];
      10'h01d: data = 32'h0c100028; // 00400074: JAL, PC<=0x00100028*4(=0x004000a0); REG[31]<=PC+4
      10'h01e: data = 32'h00000000; // 00400078: SLL, REG[0]<=REG[0]<<0;
      10'h01f: data = 32'h24020042; // 0040007c: ADDIU, REG[2]<=REG[0]+66(=0x00000042);
      10'h020: data = 32'hafc20010; // 00400080: SW, RAM[REG[30]+16]<=REG[2];
      10'h021: data = 32'hafc00014; // 00400084: SW, RAM[REG[30]+20]<=REG[0];
      10'h022: data = 32'h03c0e821; // 00400088: ADDU, REG[29]<=REG[30]+REG[0];
      10'h023: data = 32'h8fbf0114; // 0040008c: LW, REG[31]<=RAM[REG[29]+276];
      10'h024: data = 32'h8fbe0110; // 00400090: LW, REG[30]<=RAM[REG[29]+272];
      10'h025: data = 32'h27bd0118; // 00400094: ADDIU, REG[29]<=REG[29]+280(=0x00000118);
      10'h026: data = 32'h03e00008; // 00400098: JR, PC<=REG[31];
      10'h027: data = 32'h00000000; // 0040009c: SLL, REG[0]<=REG[0]<<0;
      10'h028: data = 32'h27bdfff8; // 004000a0: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h029: data = 32'hafbe0000; // 004000a4: SW, RAM[REG[29]+0]<=REG[30];
      10'h02a: data = 32'h03a0f021; // 004000a8: ADDU, REG[30]<=REG[29]+REG[0];
      10'h02b: data = 32'hafc40008; // 004000ac: SW, RAM[REG[30]+8]<=REG[4];
      10'h02c: data = 32'h081000ea; // 004000b0: J, PC<=0x001000ea*4(=0x004003a8);
      10'h02d: data = 32'h00000000; // 004000b4: SLL, REG[0]<=REG[0]<<0;
      10'h02e: data = 32'h24020300; // 004000b8: ADDIU, REG[2]<=REG[0]+768(=0x00000300);
      10'h02f: data = 32'hac400000; // 004000bc: SW, RAM[REG[2]+0]<=REG[0];
      10'h030: data = 32'h8fc20008; // 004000c0: LW, REG[2]<=RAM[REG[30]+8];
      10'h031: data = 32'h00000000; // 004000c4: SLL, REG[0]<=REG[0]<<0;
      10'h032: data = 32'h8c420000; // 004000c8: LW, REG[2]<=RAM[REG[2]+0];
      10'h033: data = 32'h00000000; // 004000cc: SLL, REG[0]<=REG[0]<<0;
      10'h034: data = 32'h2c420041; // 004000d0: SLTIU, REG[2]<=(REG[2]<65(=0x00000041))?1:0;
      10'h035: data = 32'h14400011; // 004000d4: BNE, PC<=(REG[2] != REG[0])?PC+4+17*4:PC+4;
      10'h036: data = 32'h00000000; // 004000d8: SLL, REG[0]<=REG[0]<<0;
      10'h037: data = 32'h8fc20008; // 004000dc: LW, REG[2]<=RAM[REG[30]+8];
      10'h038: data = 32'h00000000; // 004000e0: SLL, REG[0]<=REG[0]<<0;
      10'h039: data = 32'h8c420000; // 004000e4: LW, REG[2]<=RAM[REG[2]+0];
      10'h03a: data = 32'h00000000; // 004000e8: SLL, REG[0]<=REG[0]<<0;
      10'h03b: data = 32'h2c42005b; // 004000ec: SLTIU, REG[2]<=(REG[2]<91(=0x0000005b))?1:0;
      10'h03c: data = 32'h1040000a; // 004000f0: BEQ, PC<=(REG[2] == REG[0])?PC+4+10*4:PC+4;
      10'h03d: data = 32'h00000000; // 004000f4: SLL, REG[0]<=REG[0]<<0;
      10'h03e: data = 32'h24030304; // 004000f8: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h03f: data = 32'h8fc20008; // 004000fc: LW, REG[2]<=RAM[REG[30]+8];
      10'h040: data = 32'h00000000; // 00400100: SLL, REG[0]<=REG[0]<<0;
      10'h041: data = 32'h8c420000; // 00400104: LW, REG[2]<=RAM[REG[2]+0];
      10'h042: data = 32'h00000000; // 00400108: SLL, REG[0]<=REG[0]<<0;
      10'h043: data = 32'h2442ffc0; // 0040010c: ADDIU, REG[2]<=REG[2]+65472(=0x0000ffc0);
      10'h044: data = 32'hac620000; // 00400110: SW, RAM[REG[3]+0]<=REG[2];
      10'h045: data = 32'h081000e3; // 00400114: J, PC<=0x001000e3*4(=0x0040038c);
      10'h046: data = 32'h00000000; // 00400118: SLL, REG[0]<=REG[0]<<0;
      10'h047: data = 32'h8fc20008; // 0040011c: LW, REG[2]<=RAM[REG[30]+8];
      10'h048: data = 32'h00000000; // 00400120: SLL, REG[0]<=REG[0]<<0;
      10'h049: data = 32'h8c420000; // 00400124: LW, REG[2]<=RAM[REG[2]+0];
      10'h04a: data = 32'h00000000; // 00400128: SLL, REG[0]<=REG[0]<<0;
      10'h04b: data = 32'h2c420061; // 0040012c: SLTIU, REG[2]<=(REG[2]<97(=0x00000061))?1:0;
      10'h04c: data = 32'h14400011; // 00400130: BNE, PC<=(REG[2] != REG[0])?PC+4+17*4:PC+4;
      10'h04d: data = 32'h00000000; // 00400134: SLL, REG[0]<=REG[0]<<0;
      10'h04e: data = 32'h8fc20008; // 00400138: LW, REG[2]<=RAM[REG[30]+8];
      10'h04f: data = 32'h00000000; // 0040013c: SLL, REG[0]<=REG[0]<<0;
      10'h050: data = 32'h8c420000; // 00400140: LW, REG[2]<=RAM[REG[2]+0];
      10'h051: data = 32'h00000000; // 00400144: SLL, REG[0]<=REG[0]<<0;
      10'h052: data = 32'h2c42007b; // 00400148: SLTIU, REG[2]<=(REG[2]<123(=0x0000007b))?1:0;
      10'h053: data = 32'h1040000a; // 0040014c: BEQ, PC<=(REG[2] == REG[0])?PC+4+10*4:PC+4;
      10'h054: data = 32'h00000000; // 00400150: SLL, REG[0]<=REG[0]<<0;
      10'h055: data = 32'h24030304; // 00400154: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h056: data = 32'h8fc20008; // 00400158: LW, REG[2]<=RAM[REG[30]+8];
      10'h057: data = 32'h00000000; // 0040015c: SLL, REG[0]<=REG[0]<<0;
      10'h058: data = 32'h8c420000; // 00400160: LW, REG[2]<=RAM[REG[2]+0];
      10'h059: data = 32'h00000000; // 00400164: SLL, REG[0]<=REG[0]<<0;
      10'h05a: data = 32'h2442ffa0; // 00400168: ADDIU, REG[2]<=REG[2]+65440(=0x0000ffa0);
      10'h05b: data = 32'hac620000; // 0040016c: SW, RAM[REG[3]+0]<=REG[2];
      10'h05c: data = 32'h081000e3; // 00400170: J, PC<=0x001000e3*4(=0x0040038c);
      10'h05d: data = 32'h00000000; // 00400174: SLL, REG[0]<=REG[0]<<0;
      10'h05e: data = 32'h8fc20008; // 00400178: LW, REG[2]<=RAM[REG[30]+8];
      10'h05f: data = 32'h00000000; // 0040017c: SLL, REG[0]<=REG[0]<<0;
      10'h060: data = 32'h8c420000; // 00400180: LW, REG[2]<=RAM[REG[2]+0];
      10'h061: data = 32'h00000000; // 00400184: SLL, REG[0]<=REG[0]<<0;
      10'h062: data = 32'h2c420030; // 00400188: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h063: data = 32'h14400010; // 0040018c: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h064: data = 32'h00000000; // 00400190: SLL, REG[0]<=REG[0]<<0;
      10'h065: data = 32'h8fc20008; // 00400194: LW, REG[2]<=RAM[REG[30]+8];
      10'h066: data = 32'h00000000; // 00400198: SLL, REG[0]<=REG[0]<<0;
      10'h067: data = 32'h8c420000; // 0040019c: LW, REG[2]<=RAM[REG[2]+0];
      10'h068: data = 32'h00000000; // 004001a0: SLL, REG[0]<=REG[0]<<0;
      10'h069: data = 32'h2c42003a; // 004001a4: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h06a: data = 32'h10400009; // 004001a8: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h06b: data = 32'h00000000; // 004001ac: SLL, REG[0]<=REG[0]<<0;
      10'h06c: data = 32'h24020304; // 004001b0: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h06d: data = 32'h8fc30008; // 004001b4: LW, REG[3]<=RAM[REG[30]+8];
      10'h06e: data = 32'h00000000; // 004001b8: SLL, REG[0]<=REG[0]<<0;
      10'h06f: data = 32'h8c630000; // 004001bc: LW, REG[3]<=RAM[REG[3]+0];
      10'h070: data = 32'h00000000; // 004001c0: SLL, REG[0]<=REG[0]<<0;
      10'h071: data = 32'hac430000; // 004001c4: SW, RAM[REG[2]+0]<=REG[3];
      10'h072: data = 32'h081000e3; // 004001c8: J, PC<=0x001000e3*4(=0x0040038c);
      10'h073: data = 32'h00000000; // 004001cc: SLL, REG[0]<=REG[0]<<0;
      10'h074: data = 32'h8fc20008; // 004001d0: LW, REG[2]<=RAM[REG[30]+8];
      10'h075: data = 32'h00000000; // 004001d4: SLL, REG[0]<=REG[0]<<0;
      10'h076: data = 32'h8c430000; // 004001d8: LW, REG[3]<=RAM[REG[2]+0];
      10'h077: data = 32'h24020040; // 004001dc: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h078: data = 32'h14620005; // 004001e0: BNE, PC<=(REG[3] != REG[2])?PC+4+5*4:PC+4;
      10'h079: data = 32'h00000000; // 004001e4: SLL, REG[0]<=REG[0]<<0;
      10'h07a: data = 32'h24020304; // 004001e8: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h07b: data = 32'hac400000; // 004001ec: SW, RAM[REG[2]+0]<=REG[0];
      10'h07c: data = 32'h081000e3; // 004001f0: J, PC<=0x001000e3*4(=0x0040038c);
      10'h07d: data = 32'h00000000; // 004001f4: SLL, REG[0]<=REG[0]<<0;
      10'h07e: data = 32'h8fc20008; // 004001f8: LW, REG[2]<=RAM[REG[30]+8];
      10'h07f: data = 32'h00000000; // 004001fc: SLL, REG[0]<=REG[0]<<0;
      10'h080: data = 32'h8c430000; // 00400200: LW, REG[3]<=RAM[REG[2]+0];
      10'h081: data = 32'h2402005b; // 00400204: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h082: data = 32'h14620006; // 00400208: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h083: data = 32'h00000000; // 0040020c: SLL, REG[0]<=REG[0]<<0;
      10'h084: data = 32'h24030304; // 00400210: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h085: data = 32'h2402001b; // 00400214: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h086: data = 32'hac620000; // 00400218: SW, RAM[REG[3]+0]<=REG[2];
      10'h087: data = 32'h081000e3; // 0040021c: J, PC<=0x001000e3*4(=0x0040038c);
      10'h088: data = 32'h00000000; // 00400220: SLL, REG[0]<=REG[0]<<0;
      10'h089: data = 32'h8fc20008; // 00400224: LW, REG[2]<=RAM[REG[30]+8];
      10'h08a: data = 32'h00000000; // 00400228: SLL, REG[0]<=REG[0]<<0;
      10'h08b: data = 32'h8c430000; // 0040022c: LW, REG[3]<=RAM[REG[2]+0];
      10'h08c: data = 32'h2402005d; // 00400230: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h08d: data = 32'h14620006; // 00400234: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h08e: data = 32'h00000000; // 00400238: SLL, REG[0]<=REG[0]<<0;
      10'h08f: data = 32'h24030304; // 0040023c: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h090: data = 32'h2402001d; // 00400240: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h091: data = 32'hac620000; // 00400244: SW, RAM[REG[3]+0]<=REG[2];
      10'h092: data = 32'h081000e3; // 00400248: J, PC<=0x001000e3*4(=0x0040038c);
      10'h093: data = 32'h00000000; // 0040024c: SLL, REG[0]<=REG[0]<<0;
      10'h094: data = 32'h8fc20008; // 00400250: LW, REG[2]<=RAM[REG[30]+8];
      10'h095: data = 32'h00000000; // 00400254: SLL, REG[0]<=REG[0]<<0;
      10'h096: data = 32'h8c420000; // 00400258: LW, REG[2]<=RAM[REG[2]+0];
      10'h097: data = 32'h00000000; // 0040025c: SLL, REG[0]<=REG[0]<<0;
      10'h098: data = 32'h2c420020; // 00400260: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h099: data = 32'h14400010; // 00400264: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h09a: data = 32'h00000000; // 00400268: SLL, REG[0]<=REG[0]<<0;
      10'h09b: data = 32'h8fc20008; // 0040026c: LW, REG[2]<=RAM[REG[30]+8];
      10'h09c: data = 32'h00000000; // 00400270: SLL, REG[0]<=REG[0]<<0;
      10'h09d: data = 32'h8c420000; // 00400274: LW, REG[2]<=RAM[REG[2]+0];
      10'h09e: data = 32'h00000000; // 00400278: SLL, REG[0]<=REG[0]<<0;
      10'h09f: data = 32'h2c420030; // 0040027c: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h0a0: data = 32'h10400009; // 00400280: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h0a1: data = 32'h00000000; // 00400284: SLL, REG[0]<=REG[0]<<0;
      10'h0a2: data = 32'h24020304; // 00400288: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h0a3: data = 32'h8fc30008; // 0040028c: LW, REG[3]<=RAM[REG[30]+8];
      10'h0a4: data = 32'h00000000; // 00400290: SLL, REG[0]<=REG[0]<<0;
      10'h0a5: data = 32'h8c630000; // 00400294: LW, REG[3]<=RAM[REG[3]+0];
      10'h0a6: data = 32'h00000000; // 00400298: SLL, REG[0]<=REG[0]<<0;
      10'h0a7: data = 32'hac430000; // 0040029c: SW, RAM[REG[2]+0]<=REG[3];
      10'h0a8: data = 32'h081000e3; // 004002a0: J, PC<=0x001000e3*4(=0x0040038c);
      10'h0a9: data = 32'h00000000; // 004002a4: SLL, REG[0]<=REG[0]<<0;
      10'h0aa: data = 32'h8fc20008; // 004002a8: LW, REG[2]<=RAM[REG[30]+8];
      10'h0ab: data = 32'h00000000; // 004002ac: SLL, REG[0]<=REG[0]<<0;
      10'h0ac: data = 32'h8c430000; // 004002b0: LW, REG[3]<=RAM[REG[2]+0];
      10'h0ad: data = 32'h2402003f; // 004002b4: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h0ae: data = 32'h14620006; // 004002b8: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0af: data = 32'h00000000; // 004002bc: SLL, REG[0]<=REG[0]<<0;
      10'h0b0: data = 32'h24030304; // 004002c0: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h0b1: data = 32'h2402003a; // 004002c4: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h0b2: data = 32'hac620000; // 004002c8: SW, RAM[REG[3]+0]<=REG[2];
      10'h0b3: data = 32'h081000e3; // 004002cc: J, PC<=0x001000e3*4(=0x0040038c);
      10'h0b4: data = 32'h00000000; // 004002d0: SLL, REG[0]<=REG[0]<<0;
      10'h0b5: data = 32'h8fc20008; // 004002d4: LW, REG[2]<=RAM[REG[30]+8];
      10'h0b6: data = 32'h00000000; // 004002d8: SLL, REG[0]<=REG[0]<<0;
      10'h0b7: data = 32'h8c430000; // 004002dc: LW, REG[3]<=RAM[REG[2]+0];
      10'h0b8: data = 32'h2402003d; // 004002e0: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h0b9: data = 32'h14620006; // 004002e4: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0ba: data = 32'h00000000; // 004002e8: SLL, REG[0]<=REG[0]<<0;
      10'h0bb: data = 32'h24030304; // 004002ec: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h0bc: data = 32'h2402003b; // 004002f0: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h0bd: data = 32'hac620000; // 004002f4: SW, RAM[REG[3]+0]<=REG[2];
      10'h0be: data = 32'h081000e3; // 004002f8: J, PC<=0x001000e3*4(=0x0040038c);
      10'h0bf: data = 32'h00000000; // 004002fc: SLL, REG[0]<=REG[0]<<0;
      10'h0c0: data = 32'h8fc20008; // 00400300: LW, REG[2]<=RAM[REG[30]+8];
      10'h0c1: data = 32'h00000000; // 00400304: SLL, REG[0]<=REG[0]<<0;
      10'h0c2: data = 32'h8c430000; // 00400308: LW, REG[3]<=RAM[REG[2]+0];
      10'h0c3: data = 32'h2402003b; // 0040030c: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h0c4: data = 32'h14620006; // 00400310: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0c5: data = 32'h00000000; // 00400314: SLL, REG[0]<=REG[0]<<0;
      10'h0c6: data = 32'h24030304; // 00400318: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h0c7: data = 32'h2402003c; // 0040031c: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h0c8: data = 32'hac620000; // 00400320: SW, RAM[REG[3]+0]<=REG[2];
      10'h0c9: data = 32'h081000e3; // 00400324: J, PC<=0x001000e3*4(=0x0040038c);
      10'h0ca: data = 32'h00000000; // 00400328: SLL, REG[0]<=REG[0]<<0;
      10'h0cb: data = 32'h8fc20008; // 0040032c: LW, REG[2]<=RAM[REG[30]+8];
      10'h0cc: data = 32'h00000000; // 00400330: SLL, REG[0]<=REG[0]<<0;
      10'h0cd: data = 32'h8c430000; // 00400334: LW, REG[3]<=RAM[REG[2]+0];
      10'h0ce: data = 32'h2402003a; // 00400338: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h0cf: data = 32'h14620006; // 0040033c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0d0: data = 32'h00000000; // 00400340: SLL, REG[0]<=REG[0]<<0;
      10'h0d1: data = 32'h24030304; // 00400344: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h0d2: data = 32'h2402003d; // 00400348: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h0d3: data = 32'hac620000; // 0040034c: SW, RAM[REG[3]+0]<=REG[2];
      10'h0d4: data = 32'h081000e3; // 00400350: J, PC<=0x001000e3*4(=0x0040038c);
      10'h0d5: data = 32'h00000000; // 00400354: SLL, REG[0]<=REG[0]<<0;
      10'h0d6: data = 32'h8fc20008; // 00400358: LW, REG[2]<=RAM[REG[30]+8];
      10'h0d7: data = 32'h00000000; // 0040035c: SLL, REG[0]<=REG[0]<<0;
      10'h0d8: data = 32'h8c430000; // 00400360: LW, REG[3]<=RAM[REG[2]+0];
      10'h0d9: data = 32'h2402000a; // 00400364: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h0da: data = 32'h14620006; // 00400368: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0db: data = 32'h00000000; // 0040036c: SLL, REG[0]<=REG[0]<<0;
      10'h0dc: data = 32'h24030304; // 00400370: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h0dd: data = 32'h2402003e; // 00400374: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h0de: data = 32'hac620000; // 00400378: SW, RAM[REG[3]+0]<=REG[2];
      10'h0df: data = 32'h081000e3; // 0040037c: J, PC<=0x001000e3*4(=0x0040038c);
      10'h0e0: data = 32'h00000000; // 00400380: SLL, REG[0]<=REG[0]<<0;
      10'h0e1: data = 32'h24020304; // 00400384: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h0e2: data = 32'hac400000; // 00400388: SW, RAM[REG[2]+0]<=REG[0];
      10'h0e3: data = 32'h24030300; // 0040038c: ADDIU, REG[3]<=REG[0]+768(=0x00000300);
      10'h0e4: data = 32'h24020001; // 00400390: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0e5: data = 32'hac620000; // 00400394: SW, RAM[REG[3]+0]<=REG[2];
      10'h0e6: data = 32'h8fc20008; // 00400398: LW, REG[2]<=RAM[REG[30]+8];
      10'h0e7: data = 32'h00000000; // 0040039c: SLL, REG[0]<=REG[0]<<0;
      10'h0e8: data = 32'h24420004; // 004003a0: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h0e9: data = 32'hafc20008; // 004003a4: SW, RAM[REG[30]+8]<=REG[2];
      10'h0ea: data = 32'h8fc20008; // 004003a8: LW, REG[2]<=RAM[REG[30]+8];
      10'h0eb: data = 32'h00000000; // 004003ac: SLL, REG[0]<=REG[0]<<0;
      10'h0ec: data = 32'h8c420000; // 004003b0: LW, REG[2]<=RAM[REG[2]+0];
      10'h0ed: data = 32'h00000000; // 004003b4: SLL, REG[0]<=REG[0]<<0;
      10'h0ee: data = 32'h1440ff3f; // 004003b8: BNE, PC<=(REG[2] != REG[0])?PC+4+65343*4:PC+4;
      10'h0ef: data = 32'h00000000; // 004003bc: SLL, REG[0]<=REG[0]<<0;
      10'h0f0: data = 32'h03c0e821; // 004003c0: ADDU, REG[29]<=REG[30]+REG[0];
      10'h0f1: data = 32'h8fbe0000; // 004003c4: LW, REG[30]<=RAM[REG[29]+0];
      10'h0f2: data = 32'h27bd0008; // 004003c8: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h0f3: data = 32'h03e00008; // 004003cc: JR, PC<=REG[31];
      10'h0f4: data = 32'h00000000; // 004003d0: SLL, REG[0]<=REG[0]<<0;
      10'h0f5: data = 32'h00000000; // 004003d4: SLL, REG[0]<=REG[0]<<0;
      10'h0f6: data = 32'h00000000; // 004003d8: SLL, REG[0]<=REG[0]<<0;
      10'h0f7: data = 32'h00000000; // 004003dc: SLL, REG[0]<=REG[0]<<0;
    endcase
  end

  assign rom_data = data;
endmodule
