/*******************/
/* rom8x1024_sim.v */
/*******************/

//                  +----+
//  rom_addr[11:0]->|    |->rom_data[31:0]
//                  +----+

//
// ROM�ε��ҡ��������ߥ�졼������ѡ�
//

module rom8x1024_sim (rom_addr, rom_data);

  input   [11:0]  rom_addr;  // 12-bit ���ɥ쥹���ϥݡ���
  output  [31:0]  rom_data;  // 32-bit �ǡ������ϥݡ���

  reg     [31:0]  data;

  // Wire
  wire     [9:0]  word_addr; // 10-bit address, word

  assign word_addr = rom_addr[9:2];
   
  always @(word_addr) begin
    case (word_addr)
      10'h000: data = 32'he000001c; // 00400000: other type! opcode=56(10)
      10'h001: data = 32'h00000000; // 00400004: SLL, REG[0]<=REG[0]<<0;
      10'h002: data = 32'h00000000; // 00400008: SLL, REG[0]<=REG[0]<<0;
      10'h003: data = 32'h00000000; // 0040000c: SLL, REG[0]<=REG[0]<<0;
      10'h004: data = 32'h00000000; // 00400010: SLL, REG[0]<=REG[0]<<0;
      10'h005: data = 32'h00408c50; // 00400014: R type, unknown. func=16(10)
      10'h006: data = 32'h00000000; // 00400018: SLL, REG[0]<=REG[0]<<0;
      10'h007: data = 32'h00000000; // 0040001c: SLL, REG[0]<=REG[0]<<0;
      10'h008: data = 32'h27bdff60; // 00400020: ADDIU, REG[29]<=REG[29]+65376(=0x0000ff60);
      10'h009: data = 32'hafbf009c; // 00400024: SW, RAM[REG[29]+156]<=REG[31];
      10'h00a: data = 32'hafbe0098; // 00400028: SW, RAM[REG[29]+152]<=REG[30];
      10'h00b: data = 32'h03a0f021; // 0040002c: ADDU, REG[30]<=REG[29]+REG[0];
      10'h00c: data = 32'h24020048; // 00400030: ADDIU, REG[2]<=REG[0]+72(=0x00000048);
      10'h00d: data = 32'hafc20018; // 00400034: SW, RAM[REG[30]+24]<=REG[2];
      10'h00e: data = 32'h24020045; // 00400038: ADDIU, REG[2]<=REG[0]+69(=0x00000045);
      10'h00f: data = 32'hafc2001c; // 0040003c: SW, RAM[REG[30]+28]<=REG[2];
      10'h010: data = 32'h2402004c; // 00400040: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h011: data = 32'hafc20020; // 00400044: SW, RAM[REG[30]+32]<=REG[2];
      10'h012: data = 32'h2402004c; // 00400048: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h013: data = 32'hafc20024; // 0040004c: SW, RAM[REG[30]+36]<=REG[2];
      10'h014: data = 32'h2402004f; // 00400050: ADDIU, REG[2]<=REG[0]+79(=0x0000004f);
      10'h015: data = 32'hafc20028; // 00400054: SW, RAM[REG[30]+40]<=REG[2];
      10'h016: data = 32'h2402000a; // 00400058: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h017: data = 32'hafc2002c; // 0040005c: SW, RAM[REG[30]+44]<=REG[2];
      10'h018: data = 32'hafc00030; // 00400060: SW, RAM[REG[30]+48]<=REG[0];
      10'h019: data = 32'h27c20018; // 00400064: ADDIU, REG[2]<=REG[30]+24(=0x00000018);
      10'h01a: data = 32'h00402021; // 00400068: ADDU, REG[4]<=REG[2]+REG[0];
      10'h01b: data = 32'h0c100248; // 0040006c: JAL, PC<=0x00100248*4(=0x00400920); REG[31]<=PC+4
      10'h01c: data = 32'h00000000; // 00400070: SLL, REG[0]<=REG[0]<<0;
      10'h01d: data = 32'h2402004e; // 00400074: ADDIU, REG[2]<=REG[0]+78(=0x0000004e);
      10'h01e: data = 32'hafc20018; // 00400078: SW, RAM[REG[30]+24]<=REG[2];
      10'h01f: data = 32'h24020055; // 0040007c: ADDIU, REG[2]<=REG[0]+85(=0x00000055);
      10'h020: data = 32'hafc2001c; // 00400080: SW, RAM[REG[30]+28]<=REG[2];
      10'h021: data = 32'h2402004d; // 00400084: ADDIU, REG[2]<=REG[0]+77(=0x0000004d);
      10'h022: data = 32'hafc20020; // 00400088: SW, RAM[REG[30]+32]<=REG[2];
      10'h023: data = 32'h2402003d; // 0040008c: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h024: data = 32'hafc20024; // 00400090: SW, RAM[REG[30]+36]<=REG[2];
      10'h025: data = 32'hafc00028; // 00400094: SW, RAM[REG[30]+40]<=REG[0];
      10'h026: data = 32'h27c20018; // 00400098: ADDIU, REG[2]<=REG[30]+24(=0x00000018);
      10'h027: data = 32'h00402021; // 0040009c: ADDU, REG[4]<=REG[2]+REG[0];
      10'h028: data = 32'h0c100248; // 004000a0: JAL, PC<=0x00100248*4(=0x00400920); REG[31]<=PC+4
      10'h029: data = 32'h00000000; // 004000a4: SLL, REG[0]<=REG[0]<<0;
      10'h02a: data = 32'h27c20058; // 004000a8: ADDIU, REG[2]<=REG[30]+88(=0x00000058);
      10'h02b: data = 32'h00402021; // 004000ac: ADDU, REG[4]<=REG[2]+REG[0];
      10'h02c: data = 32'h0c100166; // 004000b0: JAL, PC<=0x00100166*4(=0x00400598); REG[31]<=PC+4
      10'h02d: data = 32'h00000000; // 004000b4: SLL, REG[0]<=REG[0]<<0;
      10'h02e: data = 32'h24020045; // 004000b8: ADDIU, REG[2]<=REG[0]+69(=0x00000045);
      10'h02f: data = 32'hafc20018; // 004000bc: SW, RAM[REG[30]+24]<=REG[2];
      10'h030: data = 32'h24020043; // 004000c0: ADDIU, REG[2]<=REG[0]+67(=0x00000043);
      10'h031: data = 32'hafc2001c; // 004000c4: SW, RAM[REG[30]+28]<=REG[2];
      10'h032: data = 32'h24020048; // 004000c8: ADDIU, REG[2]<=REG[0]+72(=0x00000048);
      10'h033: data = 32'hafc20020; // 004000cc: SW, RAM[REG[30]+32]<=REG[2];
      10'h034: data = 32'h2402004f; // 004000d0: ADDIU, REG[2]<=REG[0]+79(=0x0000004f);
      10'h035: data = 32'hafc20024; // 004000d4: SW, RAM[REG[30]+36]<=REG[2];
      10'h036: data = 32'h24020020; // 004000d8: ADDIU, REG[2]<=REG[0]+32(=0x00000020);
      10'h037: data = 32'hafc20028; // 004000dc: SW, RAM[REG[30]+40]<=REG[2];
      10'h038: data = 32'hafc0002c; // 004000e0: SW, RAM[REG[30]+44]<=REG[0];
      10'h039: data = 32'h27c20018; // 004000e4: ADDIU, REG[2]<=REG[30]+24(=0x00000018);
      10'h03a: data = 32'h00402021; // 004000e8: ADDU, REG[4]<=REG[2]+REG[0];
      10'h03b: data = 32'h0c100248; // 004000ec: JAL, PC<=0x00100248*4(=0x00400920); REG[31]<=PC+4
      10'h03c: data = 32'h00000000; // 004000f0: SLL, REG[0]<=REG[0]<<0;
      10'h03d: data = 32'h27c20058; // 004000f4: ADDIU, REG[2]<=REG[30]+88(=0x00000058);
      10'h03e: data = 32'h00402021; // 004000f8: ADDU, REG[4]<=REG[2]+REG[0];
      10'h03f: data = 32'h0c100248; // 004000fc: JAL, PC<=0x00100248*4(=0x00400920); REG[31]<=PC+4
      10'h040: data = 32'h00000000; // 00400100: SLL, REG[0]<=REG[0]<<0;
      10'h041: data = 32'h2402000a; // 00400104: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h042: data = 32'hafc20018; // 00400108: SW, RAM[REG[30]+24]<=REG[2];
      10'h043: data = 32'hafc0001c; // 0040010c: SW, RAM[REG[30]+28]<=REG[0];
      10'h044: data = 32'h27c20018; // 00400110: ADDIU, REG[2]<=REG[30]+24(=0x00000018);
      10'h045: data = 32'h00402021; // 00400114: ADDU, REG[4]<=REG[2]+REG[0];
      10'h046: data = 32'h0c100248; // 00400118: JAL, PC<=0x00100248*4(=0x00400920); REG[31]<=PC+4
      10'h047: data = 32'h00000000; // 0040011c: SLL, REG[0]<=REG[0]<<0;
      10'h048: data = 32'h27c20058; // 00400120: ADDIU, REG[2]<=REG[30]+88(=0x00000058);
      10'h049: data = 32'h00402021; // 00400124: ADDU, REG[4]<=REG[2]+REG[0];
      10'h04a: data = 32'h0c1000a9; // 00400128: JAL, PC<=0x001000a9*4(=0x004002a4); REG[31]<=PC+4
      10'h04b: data = 32'h00000000; // 0040012c: SLL, REG[0]<=REG[0]<<0;
      10'h04c: data = 32'hafc20010; // 00400130: SW, RAM[REG[30]+16]<=REG[2];
      10'h04d: data = 32'h24020003; // 00400134: ADDIU, REG[2]<=REG[0]+3(=0x00000003);
      10'h04e: data = 32'hafc20014; // 00400138: SW, RAM[REG[30]+20]<=REG[2];
      10'h04f: data = 32'h0810005d; // 0040013c: J, PC<=0x0010005d*4(=0x00400174);
      10'h050: data = 32'h00000000; // 00400140: SLL, REG[0]<=REG[0]<<0;
      10'h051: data = 32'h8fc40014; // 00400144: LW, REG[4]<=RAM[REG[30]+20];
      10'h052: data = 32'h0c10006c; // 00400148: JAL, PC<=0x0010006c*4(=0x004001b0); REG[31]<=PC+4
      10'h053: data = 32'h00000000; // 0040014c: SLL, REG[0]<=REG[0]<<0;
      10'h054: data = 32'h10400004; // 00400150: BEQ, PC<=(REG[2] == REG[0])?PC+4+4*4:PC+4;
      10'h055: data = 32'h00000000; // 00400154: SLL, REG[0]<=REG[0]<<0;
      10'h056: data = 32'h8fc40014; // 00400158: LW, REG[4]<=RAM[REG[30]+20];
      10'h057: data = 32'h0c10013c; // 0040015c: JAL, PC<=0x0010013c*4(=0x004004f0); REG[31]<=PC+4
      10'h058: data = 32'h00000000; // 00400160: SLL, REG[0]<=REG[0]<<0;
      10'h059: data = 32'h8fc20014; // 00400164: LW, REG[2]<=RAM[REG[30]+20];
      10'h05a: data = 32'h00000000; // 00400168: SLL, REG[0]<=REG[0]<<0;
      10'h05b: data = 32'h24420001; // 0040016c: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h05c: data = 32'hafc20014; // 00400170: SW, RAM[REG[30]+20]<=REG[2];
      10'h05d: data = 32'h8fc20014; // 00400174: LW, REG[2]<=RAM[REG[30]+20];
      10'h05e: data = 32'h8fc30010; // 00400178: LW, REG[3]<=RAM[REG[30]+16];
      10'h05f: data = 32'h00000000; // 0040017c: SLL, REG[0]<=REG[0]<<0;
      10'h060: data = 32'h0062102b; // 00400180: SLTU, REG[2]<=(REG[3]<REG[2])?1:0;
      10'h061: data = 32'h1040ffef; // 00400184: BEQ, PC<=(REG[2] == REG[0])?PC+4+65519*4:PC+4;
      10'h062: data = 32'h00000000; // 00400188: SLL, REG[0]<=REG[0]<<0;
      10'h063: data = 32'h2402000a; // 0040018c: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h064: data = 32'hafc20018; // 00400190: SW, RAM[REG[30]+24]<=REG[2];
      10'h065: data = 32'hafc0001c; // 00400194: SW, RAM[REG[30]+28]<=REG[0];
      10'h066: data = 32'h27c20018; // 00400198: ADDIU, REG[2]<=REG[30]+24(=0x00000018);
      10'h067: data = 32'h00402021; // 0040019c: ADDU, REG[4]<=REG[2]+REG[0];
      10'h068: data = 32'h0c100248; // 004001a0: JAL, PC<=0x00100248*4(=0x00400920); REG[31]<=PC+4
      10'h069: data = 32'h00000000; // 004001a4: SLL, REG[0]<=REG[0]<<0;
      10'h06a: data = 32'h0810001d; // 004001a8: J, PC<=0x0010001d*4(=0x00400074);
      10'h06b: data = 32'h00000000; // 004001ac: SLL, REG[0]<=REG[0]<<0;
      10'h06c: data = 32'h27bdffe0; // 004001b0: ADDIU, REG[29]<=REG[29]+65504(=0x0000ffe0);
      10'h06d: data = 32'hafbe0018; // 004001b4: SW, RAM[REG[29]+24]<=REG[30];
      10'h06e: data = 32'h03a0f021; // 004001b8: ADDU, REG[30]<=REG[29]+REG[0];
      10'h06f: data = 32'hafc40020; // 004001bc: SW, RAM[REG[30]+32]<=REG[4];
      10'h070: data = 32'h8fc20020; // 004001c0: LW, REG[2]<=RAM[REG[30]+32];
      10'h071: data = 32'h00000000; // 004001c4: SLL, REG[0]<=REG[0]<<0;
      10'h072: data = 32'h30420001; // 004001c8: ANDI, REG[2]<=REG[2]&0x00000001;
      10'h073: data = 32'h14400004; // 004001cc: BNE, PC<=(REG[2] != REG[0])?PC+4+4*4:PC+4;
      10'h074: data = 32'h00000000; // 004001d0: SLL, REG[0]<=REG[0]<<0;
      10'h075: data = 32'hafc00010; // 004001d4: SW, RAM[REG[30]+16]<=REG[0];
      10'h076: data = 32'h081000a3; // 004001d8: J, PC<=0x001000a3*4(=0x0040028c);
      10'h077: data = 32'h00000000; // 004001dc: SLL, REG[0]<=REG[0]<<0;
      10'h078: data = 32'h24020001; // 004001e0: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h079: data = 32'hafc20004; // 004001e4: SW, RAM[REG[30]+4]<=REG[2];
      10'h07a: data = 32'h24020003; // 004001e8: ADDIU, REG[2]<=REG[0]+3(=0x00000003);
      10'h07b: data = 32'hafc20008; // 004001ec: SW, RAM[REG[30]+8]<=REG[2];
      10'h07c: data = 32'h08100098; // 004001f0: J, PC<=0x00100098*4(=0x00400260);
      10'h07d: data = 32'h00000000; // 004001f4: SLL, REG[0]<=REG[0]<<0;
      10'h07e: data = 32'h8fc20008; // 004001f8: LW, REG[2]<=RAM[REG[30]+8];
      10'h07f: data = 32'h00000000; // 004001fc: SLL, REG[0]<=REG[0]<<0;
      10'h080: data = 32'hafc20000; // 00400200: SW, RAM[REG[30]+0]<=REG[2];
      10'h081: data = 32'h0810008e; // 00400204: J, PC<=0x0010008e*4(=0x00400238);
      10'h082: data = 32'h00000000; // 00400208: SLL, REG[0]<=REG[0]<<0;
      10'h083: data = 32'h8fc30020; // 0040020c: LW, REG[3]<=RAM[REG[30]+32];
      10'h084: data = 32'h8fc20000; // 00400210: LW, REG[2]<=RAM[REG[30]+0];
      10'h085: data = 32'h00000000; // 00400214: SLL, REG[0]<=REG[0]<<0;
      10'h086: data = 32'h14620002; // 00400218: BNE, PC<=(REG[3] != REG[2])?PC+4+2*4:PC+4;
      10'h087: data = 32'h00000000; // 0040021c: SLL, REG[0]<=REG[0]<<0;
      10'h088: data = 32'hafc00004; // 00400220: SW, RAM[REG[30]+4]<=REG[0];
      10'h089: data = 32'h8fc20000; // 00400224: LW, REG[2]<=RAM[REG[30]+0];
      10'h08a: data = 32'h8fc30008; // 00400228: LW, REG[3]<=RAM[REG[30]+8];
      10'h08b: data = 32'h00000000; // 0040022c: SLL, REG[0]<=REG[0]<<0;
      10'h08c: data = 32'h00431021; // 00400230: ADDU, REG[2]<=REG[2]+REG[3];
      10'h08d: data = 32'hafc20000; // 00400234: SW, RAM[REG[30]+0]<=REG[2];
      10'h08e: data = 32'h8fc20000; // 00400238: LW, REG[2]<=RAM[REG[30]+0];
      10'h08f: data = 32'h8fc30020; // 0040023c: LW, REG[3]<=RAM[REG[30]+32];
      10'h090: data = 32'h00000000; // 00400240: SLL, REG[0]<=REG[0]<<0;
      10'h091: data = 32'h0062102b; // 00400244: SLTU, REG[2]<=(REG[3]<REG[2])?1:0;
      10'h092: data = 32'h1040fff0; // 00400248: BEQ, PC<=(REG[2] == REG[0])?PC+4+65520*4:PC+4;
      10'h093: data = 32'h00000000; // 0040024c: SLL, REG[0]<=REG[0]<<0;
      10'h094: data = 32'h8fc20008; // 00400250: LW, REG[2]<=RAM[REG[30]+8];
      10'h095: data = 32'h00000000; // 00400254: SLL, REG[0]<=REG[0]<<0;
      10'h096: data = 32'h24420002; // 00400258: ADDIU, REG[2]<=REG[2]+2(=0x00000002);
      10'h097: data = 32'hafc20008; // 0040025c: SW, RAM[REG[30]+8]<=REG[2];
      10'h098: data = 32'h8fc20020; // 00400260: LW, REG[2]<=RAM[REG[30]+32];
      10'h099: data = 32'h00000000; // 00400264: SLL, REG[0]<=REG[0]<<0;
      10'h09a: data = 32'h00021842; // 00400268: SRL, REG[3]<=REG[2]>>1;
      10'h09b: data = 32'h8fc20008; // 0040026c: LW, REG[2]<=RAM[REG[30]+8];
      10'h09c: data = 32'h00000000; // 00400270: SLL, REG[0]<=REG[0]<<0;
      10'h09d: data = 32'h0043102b; // 00400274: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h09e: data = 32'h1440ffdf; // 00400278: BNE, PC<=(REG[2] != REG[0])?PC+4+65503*4:PC+4;
      10'h09f: data = 32'h00000000; // 0040027c: SLL, REG[0]<=REG[0]<<0;
      10'h0a0: data = 32'h8fc20004; // 00400280: LW, REG[2]<=RAM[REG[30]+4];
      10'h0a1: data = 32'h00000000; // 00400284: SLL, REG[0]<=REG[0]<<0;
      10'h0a2: data = 32'hafc20010; // 00400288: SW, RAM[REG[30]+16]<=REG[2];
      10'h0a3: data = 32'h8fc20010; // 0040028c: LW, REG[2]<=RAM[REG[30]+16];
      10'h0a4: data = 32'h03c0e821; // 00400290: ADDU, REG[29]<=REG[30]+REG[0];
      10'h0a5: data = 32'h8fbe0018; // 00400294: LW, REG[30]<=RAM[REG[29]+24];
      10'h0a6: data = 32'h27bd0020; // 00400298: ADDIU, REG[29]<=REG[29]+32(=0x00000020);
      10'h0a7: data = 32'h03e00008; // 0040029c: JR, PC<=REG[31];
      10'h0a8: data = 32'h00000000; // 004002a0: SLL, REG[0]<=REG[0]<<0;
      10'h0a9: data = 32'h27bdffe8; // 004002a4: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h0aa: data = 32'hafbe0010; // 004002a8: SW, RAM[REG[29]+16]<=REG[30];
      10'h0ab: data = 32'h03a0f021; // 004002ac: ADDU, REG[30]<=REG[29]+REG[0];
      10'h0ac: data = 32'hafc40018; // 004002b0: SW, RAM[REG[30]+24]<=REG[4];
      10'h0ad: data = 32'h8fc20018; // 004002b4: LW, REG[2]<=RAM[REG[30]+24];
      10'h0ae: data = 32'h00000000; // 004002b8: SLL, REG[0]<=REG[0]<<0;
      10'h0af: data = 32'hafc20008; // 004002bc: SW, RAM[REG[30]+8]<=REG[2];
      10'h0b0: data = 32'hafc00004; // 004002c0: SW, RAM[REG[30]+4]<=REG[0];
      10'h0b1: data = 32'h081000bb; // 004002c4: J, PC<=0x001000bb*4(=0x004002ec);
      10'h0b2: data = 32'h00000000; // 004002c8: SLL, REG[0]<=REG[0]<<0;
      10'h0b3: data = 32'h8fc20008; // 004002cc: LW, REG[2]<=RAM[REG[30]+8];
      10'h0b4: data = 32'h00000000; // 004002d0: SLL, REG[0]<=REG[0]<<0;
      10'h0b5: data = 32'h24420004; // 004002d4: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h0b6: data = 32'hafc20008; // 004002d8: SW, RAM[REG[30]+8]<=REG[2];
      10'h0b7: data = 32'h8fc20004; // 004002dc: LW, REG[2]<=RAM[REG[30]+4];
      10'h0b8: data = 32'h00000000; // 004002e0: SLL, REG[0]<=REG[0]<<0;
      10'h0b9: data = 32'h24420001; // 004002e4: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h0ba: data = 32'hafc20004; // 004002e8: SW, RAM[REG[30]+4]<=REG[2];
      10'h0bb: data = 32'h8fc20008; // 004002ec: LW, REG[2]<=RAM[REG[30]+8];
      10'h0bc: data = 32'h00000000; // 004002f0: SLL, REG[0]<=REG[0]<<0;
      10'h0bd: data = 32'h8c420000; // 004002f4: LW, REG[2]<=RAM[REG[2]+0];
      10'h0be: data = 32'h00000000; // 004002f8: SLL, REG[0]<=REG[0]<<0;
      10'h0bf: data = 32'h1440fff3; // 004002fc: BNE, PC<=(REG[2] != REG[0])?PC+4+65523*4:PC+4;
      10'h0c0: data = 32'h00000000; // 00400300: SLL, REG[0]<=REG[0]<<0;
      10'h0c1: data = 32'hafc00000; // 00400304: SW, RAM[REG[30]+0]<=REG[0];
      10'h0c2: data = 32'h8fc20018; // 00400308: LW, REG[2]<=RAM[REG[30]+24];
      10'h0c3: data = 32'h00000000; // 0040030c: SLL, REG[0]<=REG[0]<<0;
      10'h0c4: data = 32'hafc20008; // 00400310: SW, RAM[REG[30]+8]<=REG[2];
      10'h0c5: data = 32'h8fc30004; // 00400314: LW, REG[3]<=RAM[REG[30]+4];
      10'h0c6: data = 32'h24020001; // 00400318: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0c7: data = 32'h14620009; // 0040031c: BNE, PC<=(REG[3] != REG[2])?PC+4+9*4:PC+4;
      10'h0c8: data = 32'h00000000; // 00400320: SLL, REG[0]<=REG[0]<<0;
      10'h0c9: data = 32'h8fc20008; // 00400324: LW, REG[2]<=RAM[REG[30]+8];
      10'h0ca: data = 32'h00000000; // 00400328: SLL, REG[0]<=REG[0]<<0;
      10'h0cb: data = 32'h8c420000; // 0040032c: LW, REG[2]<=RAM[REG[2]+0];
      10'h0cc: data = 32'h00000000; // 00400330: SLL, REG[0]<=REG[0]<<0;
      10'h0cd: data = 32'h2442ffd0; // 00400334: ADDIU, REG[2]<=REG[2]+65488(=0x0000ffd0);
      10'h0ce: data = 32'hafc20000; // 00400338: SW, RAM[REG[30]+0]<=REG[2];
      10'h0cf: data = 32'h08100136; // 0040033c: J, PC<=0x00100136*4(=0x004004d8);
      10'h0d0: data = 32'h00000000; // 00400340: SLL, REG[0]<=REG[0]<<0;
      10'h0d1: data = 32'h8fc30004; // 00400344: LW, REG[3]<=RAM[REG[30]+4];
      10'h0d2: data = 32'h24020002; // 00400348: ADDIU, REG[2]<=REG[0]+2(=0x00000002);
      10'h0d3: data = 32'h14620024; // 0040034c: BNE, PC<=(REG[3] != REG[2])?PC+4+36*4:PC+4;
      10'h0d4: data = 32'h00000000; // 00400350: SLL, REG[0]<=REG[0]<<0;
      10'h0d5: data = 32'hafc00004; // 00400354: SW, RAM[REG[30]+4]<=REG[0];
      10'h0d6: data = 32'h081000e0; // 00400358: J, PC<=0x001000e0*4(=0x00400380);
      10'h0d7: data = 32'h00000000; // 0040035c: SLL, REG[0]<=REG[0]<<0;
      10'h0d8: data = 32'h8fc20000; // 00400360: LW, REG[2]<=RAM[REG[30]+0];
      10'h0d9: data = 32'h00000000; // 00400364: SLL, REG[0]<=REG[0]<<0;
      10'h0da: data = 32'h2442000a; // 00400368: ADDIU, REG[2]<=REG[2]+10(=0x0000000a);
      10'h0db: data = 32'hafc20000; // 0040036c: SW, RAM[REG[30]+0]<=REG[2];
      10'h0dc: data = 32'h8fc20004; // 00400370: LW, REG[2]<=RAM[REG[30]+4];
      10'h0dd: data = 32'h00000000; // 00400374: SLL, REG[0]<=REG[0]<<0;
      10'h0de: data = 32'h24420001; // 00400378: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h0df: data = 32'hafc20004; // 0040037c: SW, RAM[REG[30]+4]<=REG[2];
      10'h0e0: data = 32'h8fc20008; // 00400380: LW, REG[2]<=RAM[REG[30]+8];
      10'h0e1: data = 32'h00000000; // 00400384: SLL, REG[0]<=REG[0]<<0;
      10'h0e2: data = 32'h8c420000; // 00400388: LW, REG[2]<=RAM[REG[2]+0];
      10'h0e3: data = 32'h00000000; // 0040038c: SLL, REG[0]<=REG[0]<<0;
      10'h0e4: data = 32'h2443ffd0; // 00400390: ADDIU, REG[3]<=REG[2]+65488(=0x0000ffd0);
      10'h0e5: data = 32'h8fc20004; // 00400394: LW, REG[2]<=RAM[REG[30]+4];
      10'h0e6: data = 32'h00000000; // 00400398: SLL, REG[0]<=REG[0]<<0;
      10'h0e7: data = 32'h0043102b; // 0040039c: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h0e8: data = 32'h1440ffef; // 004003a0: BNE, PC<=(REG[2] != REG[0])?PC+4+65519*4:PC+4;
      10'h0e9: data = 32'h00000000; // 004003a4: SLL, REG[0]<=REG[0]<<0;
      10'h0ea: data = 32'h8fc20008; // 004003a8: LW, REG[2]<=RAM[REG[30]+8];
      10'h0eb: data = 32'h00000000; // 004003ac: SLL, REG[0]<=REG[0]<<0;
      10'h0ec: data = 32'h24420004; // 004003b0: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h0ed: data = 32'hafc20008; // 004003b4: SW, RAM[REG[30]+8]<=REG[2];
      10'h0ee: data = 32'h8fc20008; // 004003b8: LW, REG[2]<=RAM[REG[30]+8];
      10'h0ef: data = 32'h00000000; // 004003bc: SLL, REG[0]<=REG[0]<<0;
      10'h0f0: data = 32'h8c430000; // 004003c0: LW, REG[3]<=RAM[REG[2]+0];
      10'h0f1: data = 32'h8fc20000; // 004003c4: LW, REG[2]<=RAM[REG[30]+0];
      10'h0f2: data = 32'h00000000; // 004003c8: SLL, REG[0]<=REG[0]<<0;
      10'h0f3: data = 32'h00621021; // 004003cc: ADDU, REG[2]<=REG[3]+REG[2];
      10'h0f4: data = 32'h2442ffd0; // 004003d0: ADDIU, REG[2]<=REG[2]+65488(=0x0000ffd0);
      10'h0f5: data = 32'hafc20000; // 004003d4: SW, RAM[REG[30]+0]<=REG[2];
      10'h0f6: data = 32'h08100136; // 004003d8: J, PC<=0x00100136*4(=0x004004d8);
      10'h0f7: data = 32'h00000000; // 004003dc: SLL, REG[0]<=REG[0]<<0;
      10'h0f8: data = 32'h8fc30004; // 004003e0: LW, REG[3]<=RAM[REG[30]+4];
      10'h0f9: data = 32'h24020003; // 004003e4: ADDIU, REG[2]<=REG[0]+3(=0x00000003);
      10'h0fa: data = 32'h1462003b; // 004003e8: BNE, PC<=(REG[3] != REG[2])?PC+4+59*4:PC+4;
      10'h0fb: data = 32'h00000000; // 004003ec: SLL, REG[0]<=REG[0]<<0;
      10'h0fc: data = 32'hafc00004; // 004003f0: SW, RAM[REG[30]+4]<=REG[0];
      10'h0fd: data = 32'h08100107; // 004003f4: J, PC<=0x00100107*4(=0x0040041c);
      10'h0fe: data = 32'h00000000; // 004003f8: SLL, REG[0]<=REG[0]<<0;
      10'h0ff: data = 32'h8fc20000; // 004003fc: LW, REG[2]<=RAM[REG[30]+0];
      10'h100: data = 32'h00000000; // 00400400: SLL, REG[0]<=REG[0]<<0;
      10'h101: data = 32'h24420064; // 00400404: ADDIU, REG[2]<=REG[2]+100(=0x00000064);
      10'h102: data = 32'hafc20000; // 00400408: SW, RAM[REG[30]+0]<=REG[2];
      10'h103: data = 32'h8fc20004; // 0040040c: LW, REG[2]<=RAM[REG[30]+4];
      10'h104: data = 32'h00000000; // 00400410: SLL, REG[0]<=REG[0]<<0;
      10'h105: data = 32'h24420001; // 00400414: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h106: data = 32'hafc20004; // 00400418: SW, RAM[REG[30]+4]<=REG[2];
      10'h107: data = 32'h8fc20008; // 0040041c: LW, REG[2]<=RAM[REG[30]+8];
      10'h108: data = 32'h00000000; // 00400420: SLL, REG[0]<=REG[0]<<0;
      10'h109: data = 32'h8c420000; // 00400424: LW, REG[2]<=RAM[REG[2]+0];
      10'h10a: data = 32'h00000000; // 00400428: SLL, REG[0]<=REG[0]<<0;
      10'h10b: data = 32'h2443ffd0; // 0040042c: ADDIU, REG[3]<=REG[2]+65488(=0x0000ffd0);
      10'h10c: data = 32'h8fc20004; // 00400430: LW, REG[2]<=RAM[REG[30]+4];
      10'h10d: data = 32'h00000000; // 00400434: SLL, REG[0]<=REG[0]<<0;
      10'h10e: data = 32'h0043102b; // 00400438: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h10f: data = 32'h1440ffef; // 0040043c: BNE, PC<=(REG[2] != REG[0])?PC+4+65519*4:PC+4;
      10'h110: data = 32'h00000000; // 00400440: SLL, REG[0]<=REG[0]<<0;
      10'h111: data = 32'h8fc20008; // 00400444: LW, REG[2]<=RAM[REG[30]+8];
      10'h112: data = 32'h00000000; // 00400448: SLL, REG[0]<=REG[0]<<0;
      10'h113: data = 32'h24420004; // 0040044c: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h114: data = 32'hafc20008; // 00400450: SW, RAM[REG[30]+8]<=REG[2];
      10'h115: data = 32'hafc00004; // 00400454: SW, RAM[REG[30]+4]<=REG[0];
      10'h116: data = 32'h08100120; // 00400458: J, PC<=0x00100120*4(=0x00400480);
      10'h117: data = 32'h00000000; // 0040045c: SLL, REG[0]<=REG[0]<<0;
      10'h118: data = 32'h8fc20000; // 00400460: LW, REG[2]<=RAM[REG[30]+0];
      10'h119: data = 32'h00000000; // 00400464: SLL, REG[0]<=REG[0]<<0;
      10'h11a: data = 32'h2442000a; // 00400468: ADDIU, REG[2]<=REG[2]+10(=0x0000000a);
      10'h11b: data = 32'hafc20000; // 0040046c: SW, RAM[REG[30]+0]<=REG[2];
      10'h11c: data = 32'h8fc20004; // 00400470: LW, REG[2]<=RAM[REG[30]+4];
      10'h11d: data = 32'h00000000; // 00400474: SLL, REG[0]<=REG[0]<<0;
      10'h11e: data = 32'h24420001; // 00400478: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h11f: data = 32'hafc20004; // 0040047c: SW, RAM[REG[30]+4]<=REG[2];
      10'h120: data = 32'h8fc20008; // 00400480: LW, REG[2]<=RAM[REG[30]+8];
      10'h121: data = 32'h00000000; // 00400484: SLL, REG[0]<=REG[0]<<0;
      10'h122: data = 32'h8c420000; // 00400488: LW, REG[2]<=RAM[REG[2]+0];
      10'h123: data = 32'h00000000; // 0040048c: SLL, REG[0]<=REG[0]<<0;
      10'h124: data = 32'h2443ffd0; // 00400490: ADDIU, REG[3]<=REG[2]+65488(=0x0000ffd0);
      10'h125: data = 32'h8fc20004; // 00400494: LW, REG[2]<=RAM[REG[30]+4];
      10'h126: data = 32'h00000000; // 00400498: SLL, REG[0]<=REG[0]<<0;
      10'h127: data = 32'h0043102b; // 0040049c: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h128: data = 32'h1440ffef; // 004004a0: BNE, PC<=(REG[2] != REG[0])?PC+4+65519*4:PC+4;
      10'h129: data = 32'h00000000; // 004004a4: SLL, REG[0]<=REG[0]<<0;
      10'h12a: data = 32'h8fc20008; // 004004a8: LW, REG[2]<=RAM[REG[30]+8];
      10'h12b: data = 32'h00000000; // 004004ac: SLL, REG[0]<=REG[0]<<0;
      10'h12c: data = 32'h24420004; // 004004b0: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h12d: data = 32'hafc20008; // 004004b4: SW, RAM[REG[30]+8]<=REG[2];
      10'h12e: data = 32'h8fc20008; // 004004b8: LW, REG[2]<=RAM[REG[30]+8];
      10'h12f: data = 32'h00000000; // 004004bc: SLL, REG[0]<=REG[0]<<0;
      10'h130: data = 32'h8c430000; // 004004c0: LW, REG[3]<=RAM[REG[2]+0];
      10'h131: data = 32'h8fc20000; // 004004c4: LW, REG[2]<=RAM[REG[30]+0];
      10'h132: data = 32'h00000000; // 004004c8: SLL, REG[0]<=REG[0]<<0;
      10'h133: data = 32'h00621021; // 004004cc: ADDU, REG[2]<=REG[3]+REG[2];
      10'h134: data = 32'h2442ffd0; // 004004d0: ADDIU, REG[2]<=REG[2]+65488(=0x0000ffd0);
      10'h135: data = 32'hafc20000; // 004004d4: SW, RAM[REG[30]+0]<=REG[2];
      10'h136: data = 32'h8fc20000; // 004004d8: LW, REG[2]<=RAM[REG[30]+0];
      10'h137: data = 32'h03c0e821; // 004004dc: ADDU, REG[29]<=REG[30]+REG[0];
      10'h138: data = 32'h8fbe0010; // 004004e0: LW, REG[30]<=RAM[REG[29]+16];
      10'h139: data = 32'h27bd0018; // 004004e4: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h13a: data = 32'h03e00008; // 004004e8: JR, PC<=REG[31];
      10'h13b: data = 32'h00000000; // 004004ec: SLL, REG[0]<=REG[0]<<0;
      10'h13c: data = 32'h27bdffd0; // 004004f0: ADDIU, REG[29]<=REG[29]+65488(=0x0000ffd0);
      10'h13d: data = 32'hafbf002c; // 004004f4: SW, RAM[REG[29]+44]<=REG[31];
      10'h13e: data = 32'hafbe0028; // 004004f8: SW, RAM[REG[29]+40]<=REG[30];
      10'h13f: data = 32'h03a0f021; // 004004fc: ADDU, REG[30]<=REG[29]+REG[0];
      10'h140: data = 32'hafc40030; // 00400500: SW, RAM[REG[30]+48]<=REG[4];
      10'h141: data = 32'hafc00010; // 00400504: SW, RAM[REG[30]+16]<=REG[0];
      10'h142: data = 32'h0810014c; // 00400508: J, PC<=0x0010014c*4(=0x00400530);
      10'h143: data = 32'h00000000; // 0040050c: SLL, REG[0]<=REG[0]<<0;
      10'h144: data = 32'h8fc20030; // 00400510: LW, REG[2]<=RAM[REG[30]+48];
      10'h145: data = 32'h00000000; // 00400514: SLL, REG[0]<=REG[0]<<0;
      10'h146: data = 32'h2442fff6; // 00400518: ADDIU, REG[2]<=REG[2]+65526(=0x0000fff6);
      10'h147: data = 32'hafc20030; // 0040051c: SW, RAM[REG[30]+48]<=REG[2];
      10'h148: data = 32'h8fc20010; // 00400520: LW, REG[2]<=RAM[REG[30]+16];
      10'h149: data = 32'h00000000; // 00400524: SLL, REG[0]<=REG[0]<<0;
      10'h14a: data = 32'h24420001; // 00400528: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h14b: data = 32'hafc20010; // 0040052c: SW, RAM[REG[30]+16]<=REG[2];
      10'h14c: data = 32'h8fc20030; // 00400530: LW, REG[2]<=RAM[REG[30]+48];
      10'h14d: data = 32'h00000000; // 00400534: SLL, REG[0]<=REG[0]<<0;
      10'h14e: data = 32'h2c42000a; // 00400538: SLTIU, REG[2]<=(REG[2]<10(=0x0000000a))?1:0;
      10'h14f: data = 32'h1040fff4; // 0040053c: BEQ, PC<=(REG[2] == REG[0])?PC+4+65524*4:PC+4;
      10'h150: data = 32'h00000000; // 00400540: SLL, REG[0]<=REG[0]<<0;
      10'h151: data = 32'h8fc20010; // 00400544: LW, REG[2]<=RAM[REG[30]+16];
      10'h152: data = 32'h00000000; // 00400548: SLL, REG[0]<=REG[0]<<0;
      10'h153: data = 32'h24420030; // 0040054c: ADDIU, REG[2]<=REG[2]+48(=0x00000030);
      10'h154: data = 32'hafc20014; // 00400550: SW, RAM[REG[30]+20]<=REG[2];
      10'h155: data = 32'h8fc20030; // 00400554: LW, REG[2]<=RAM[REG[30]+48];
      10'h156: data = 32'h00000000; // 00400558: SLL, REG[0]<=REG[0]<<0;
      10'h157: data = 32'h24420030; // 0040055c: ADDIU, REG[2]<=REG[2]+48(=0x00000030);
      10'h158: data = 32'hafc20018; // 00400560: SW, RAM[REG[30]+24]<=REG[2];
      10'h159: data = 32'h24020020; // 00400564: ADDIU, REG[2]<=REG[0]+32(=0x00000020);
      10'h15a: data = 32'hafc2001c; // 00400568: SW, RAM[REG[30]+28]<=REG[2];
      10'h15b: data = 32'hafc00020; // 0040056c: SW, RAM[REG[30]+32]<=REG[0];
      10'h15c: data = 32'h27c20014; // 00400570: ADDIU, REG[2]<=REG[30]+20(=0x00000014);
      10'h15d: data = 32'h00402021; // 00400574: ADDU, REG[4]<=REG[2]+REG[0];
      10'h15e: data = 32'h0c100248; // 00400578: JAL, PC<=0x00100248*4(=0x00400920); REG[31]<=PC+4
      10'h15f: data = 32'h00000000; // 0040057c: SLL, REG[0]<=REG[0]<<0;
      10'h160: data = 32'h03c0e821; // 00400580: ADDU, REG[29]<=REG[30]+REG[0];
      10'h161: data = 32'h8fbf002c; // 00400584: LW, REG[31]<=RAM[REG[29]+44];
      10'h162: data = 32'h8fbe0028; // 00400588: LW, REG[30]<=RAM[REG[29]+40];
      10'h163: data = 32'h27bd0030; // 0040058c: ADDIU, REG[29]<=REG[29]+48(=0x00000030);
      10'h164: data = 32'h03e00008; // 00400590: JR, PC<=REG[31];
      10'h165: data = 32'h00000000; // 00400594: SLL, REG[0]<=REG[0]<<0;
      10'h166: data = 32'h27bdfff8; // 00400598: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h167: data = 32'hafbe0000; // 0040059c: SW, RAM[REG[29]+0]<=REG[30];
      10'h168: data = 32'h03a0f021; // 004005a0: ADDU, REG[30]<=REG[29]+REG[0];
      10'h169: data = 32'hafc40008; // 004005a4: SW, RAM[REG[30]+8]<=REG[4];
      10'h16a: data = 32'h24020308; // 004005a8: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h16b: data = 32'hac400000; // 004005ac: SW, RAM[REG[2]+0]<=REG[0];
      10'h16c: data = 32'h2403030c; // 004005b0: ADDIU, REG[3]<=REG[0]+780(=0x0000030c);
      10'h16d: data = 32'h24020001; // 004005b4: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h16e: data = 32'hac620000; // 004005b8: SW, RAM[REG[3]+0]<=REG[2];
      10'h16f: data = 32'h24030308; // 004005bc: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h170: data = 32'h24020001; // 004005c0: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h171: data = 32'hac620000; // 004005c4: SW, RAM[REG[3]+0]<=REG[2];
      10'h172: data = 32'h24020308; // 004005c8: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h173: data = 32'hac400000; // 004005cc: SW, RAM[REG[2]+0]<=REG[0];
      10'h174: data = 32'h24030308; // 004005d0: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h175: data = 32'h24020001; // 004005d4: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h176: data = 32'hac620000; // 004005d8: SW, RAM[REG[3]+0]<=REG[2];
      10'h177: data = 32'h0810017e; // 004005dc: J, PC<=0x0010017e*4(=0x004005f8);
      10'h178: data = 32'h00000000; // 004005e0: SLL, REG[0]<=REG[0]<<0;
      10'h179: data = 32'h24020308; // 004005e4: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h17a: data = 32'hac400000; // 004005e8: SW, RAM[REG[2]+0]<=REG[0];
      10'h17b: data = 32'h24030308; // 004005ec: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h17c: data = 32'h24020001; // 004005f0: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h17d: data = 32'hac620000; // 004005f4: SW, RAM[REG[3]+0]<=REG[2];
      10'h17e: data = 32'h24020310; // 004005f8: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h17f: data = 32'h8c430000; // 004005fc: LW, REG[3]<=RAM[REG[2]+0];
      10'h180: data = 32'h2402ffff; // 00400600: ADDIU, REG[2]<=REG[0]+65535(=0x0000ffff);
      10'h181: data = 32'h1062fff7; // 00400604: BEQ, PC<=(REG[3] == REG[2])?PC+4+65527*4:PC+4;
      10'h182: data = 32'h00000000; // 00400608: SLL, REG[0]<=REG[0]<<0;
      10'h183: data = 32'h0810022c; // 0040060c: J, PC<=0x0010022c*4(=0x004008b0);
      10'h184: data = 32'h00000000; // 00400610: SLL, REG[0]<=REG[0]<<0;
      10'h185: data = 32'h8fc20008; // 00400614: LW, REG[2]<=RAM[REG[30]+8];
      10'h186: data = 32'h00000000; // 00400618: SLL, REG[0]<=REG[0]<<0;
      10'h187: data = 32'h8c420000; // 0040061c: LW, REG[2]<=RAM[REG[2]+0];
      10'h188: data = 32'h00000000; // 00400620: SLL, REG[0]<=REG[0]<<0;
      10'h189: data = 32'h10400012; // 00400624: BEQ, PC<=(REG[2] == REG[0])?PC+4+18*4:PC+4;
      10'h18a: data = 32'h00000000; // 00400628: SLL, REG[0]<=REG[0]<<0;
      10'h18b: data = 32'h8fc20008; // 0040062c: LW, REG[2]<=RAM[REG[30]+8];
      10'h18c: data = 32'h00000000; // 00400630: SLL, REG[0]<=REG[0]<<0;
      10'h18d: data = 32'h8c420000; // 00400634: LW, REG[2]<=RAM[REG[2]+0];
      10'h18e: data = 32'h00000000; // 00400638: SLL, REG[0]<=REG[0]<<0;
      10'h18f: data = 32'h2c42001b; // 0040063c: SLTIU, REG[2]<=(REG[2]<27(=0x0000001b))?1:0;
      10'h190: data = 32'h1040000b; // 00400640: BEQ, PC<=(REG[2] == REG[0])?PC+4+11*4:PC+4;
      10'h191: data = 32'h00000000; // 00400644: SLL, REG[0]<=REG[0]<<0;
      10'h192: data = 32'h8fc20008; // 00400648: LW, REG[2]<=RAM[REG[30]+8];
      10'h193: data = 32'h00000000; // 0040064c: SLL, REG[0]<=REG[0]<<0;
      10'h194: data = 32'h8c420000; // 00400650: LW, REG[2]<=RAM[REG[2]+0];
      10'h195: data = 32'h00000000; // 00400654: SLL, REG[0]<=REG[0]<<0;
      10'h196: data = 32'h24430040; // 00400658: ADDIU, REG[3]<=REG[2]+64(=0x00000040);
      10'h197: data = 32'h8fc20008; // 0040065c: LW, REG[2]<=RAM[REG[30]+8];
      10'h198: data = 32'h00000000; // 00400660: SLL, REG[0]<=REG[0]<<0;
      10'h199: data = 32'hac430000; // 00400664: SW, RAM[REG[2]+0]<=REG[3];
      10'h19a: data = 32'h08100223; // 00400668: J, PC<=0x00100223*4(=0x0040088c);
      10'h19b: data = 32'h00000000; // 0040066c: SLL, REG[0]<=REG[0]<<0;
      10'h19c: data = 32'h8fc20008; // 00400670: LW, REG[2]<=RAM[REG[30]+8];
      10'h19d: data = 32'h00000000; // 00400674: SLL, REG[0]<=REG[0]<<0;
      10'h19e: data = 32'h8c420000; // 00400678: LW, REG[2]<=RAM[REG[2]+0];
      10'h19f: data = 32'h00000000; // 0040067c: SLL, REG[0]<=REG[0]<<0;
      10'h1a0: data = 32'h2c420030; // 00400680: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h1a1: data = 32'h14400010; // 00400684: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h1a2: data = 32'h00000000; // 00400688: SLL, REG[0]<=REG[0]<<0;
      10'h1a3: data = 32'h8fc20008; // 0040068c: LW, REG[2]<=RAM[REG[30]+8];
      10'h1a4: data = 32'h00000000; // 00400690: SLL, REG[0]<=REG[0]<<0;
      10'h1a5: data = 32'h8c420000; // 00400694: LW, REG[2]<=RAM[REG[2]+0];
      10'h1a6: data = 32'h00000000; // 00400698: SLL, REG[0]<=REG[0]<<0;
      10'h1a7: data = 32'h2c42003a; // 0040069c: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h1a8: data = 32'h10400009; // 004006a0: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h1a9: data = 32'h00000000; // 004006a4: SLL, REG[0]<=REG[0]<<0;
      10'h1aa: data = 32'h8fc20008; // 004006a8: LW, REG[2]<=RAM[REG[30]+8];
      10'h1ab: data = 32'h00000000; // 004006ac: SLL, REG[0]<=REG[0]<<0;
      10'h1ac: data = 32'h8c430000; // 004006b0: LW, REG[3]<=RAM[REG[2]+0];
      10'h1ad: data = 32'h8fc20008; // 004006b4: LW, REG[2]<=RAM[REG[30]+8];
      10'h1ae: data = 32'h00000000; // 004006b8: SLL, REG[0]<=REG[0]<<0;
      10'h1af: data = 32'hac430000; // 004006bc: SW, RAM[REG[2]+0]<=REG[3];
      10'h1b0: data = 32'h08100223; // 004006c0: J, PC<=0x00100223*4(=0x0040088c);
      10'h1b1: data = 32'h00000000; // 004006c4: SLL, REG[0]<=REG[0]<<0;
      10'h1b2: data = 32'h8fc20008; // 004006c8: LW, REG[2]<=RAM[REG[30]+8];
      10'h1b3: data = 32'h00000000; // 004006cc: SLL, REG[0]<=REG[0]<<0;
      10'h1b4: data = 32'h8c420000; // 004006d0: LW, REG[2]<=RAM[REG[2]+0];
      10'h1b5: data = 32'h00000000; // 004006d4: SLL, REG[0]<=REG[0]<<0;
      10'h1b6: data = 32'h14400006; // 004006d8: BNE, PC<=(REG[2] != REG[0])?PC+4+6*4:PC+4;
      10'h1b7: data = 32'h00000000; // 004006dc: SLL, REG[0]<=REG[0]<<0;
      10'h1b8: data = 32'h8fc30008; // 004006e0: LW, REG[3]<=RAM[REG[30]+8];
      10'h1b9: data = 32'h24020040; // 004006e4: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h1ba: data = 32'hac620000; // 004006e8: SW, RAM[REG[3]+0]<=REG[2];
      10'h1bb: data = 32'h08100223; // 004006ec: J, PC<=0x00100223*4(=0x0040088c);
      10'h1bc: data = 32'h00000000; // 004006f0: SLL, REG[0]<=REG[0]<<0;
      10'h1bd: data = 32'h8fc20008; // 004006f4: LW, REG[2]<=RAM[REG[30]+8];
      10'h1be: data = 32'h00000000; // 004006f8: SLL, REG[0]<=REG[0]<<0;
      10'h1bf: data = 32'h8c430000; // 004006fc: LW, REG[3]<=RAM[REG[2]+0];
      10'h1c0: data = 32'h2402001b; // 00400700: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h1c1: data = 32'h14620006; // 00400704: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1c2: data = 32'h00000000; // 00400708: SLL, REG[0]<=REG[0]<<0;
      10'h1c3: data = 32'h8fc30008; // 0040070c: LW, REG[3]<=RAM[REG[30]+8];
      10'h1c4: data = 32'h2402005b; // 00400710: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h1c5: data = 32'hac620000; // 00400714: SW, RAM[REG[3]+0]<=REG[2];
      10'h1c6: data = 32'h08100223; // 00400718: J, PC<=0x00100223*4(=0x0040088c);
      10'h1c7: data = 32'h00000000; // 0040071c: SLL, REG[0]<=REG[0]<<0;
      10'h1c8: data = 32'h8fc20008; // 00400720: LW, REG[2]<=RAM[REG[30]+8];
      10'h1c9: data = 32'h00000000; // 00400724: SLL, REG[0]<=REG[0]<<0;
      10'h1ca: data = 32'h8c430000; // 00400728: LW, REG[3]<=RAM[REG[2]+0];
      10'h1cb: data = 32'h2402001d; // 0040072c: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h1cc: data = 32'h14620006; // 00400730: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1cd: data = 32'h00000000; // 00400734: SLL, REG[0]<=REG[0]<<0;
      10'h1ce: data = 32'h8fc30008; // 00400738: LW, REG[3]<=RAM[REG[30]+8];
      10'h1cf: data = 32'h2402005d; // 0040073c: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h1d0: data = 32'hac620000; // 00400740: SW, RAM[REG[3]+0]<=REG[2];
      10'h1d1: data = 32'h08100223; // 00400744: J, PC<=0x00100223*4(=0x0040088c);
      10'h1d2: data = 32'h00000000; // 00400748: SLL, REG[0]<=REG[0]<<0;
      10'h1d3: data = 32'h8fc20008; // 0040074c: LW, REG[2]<=RAM[REG[30]+8];
      10'h1d4: data = 32'h00000000; // 00400750: SLL, REG[0]<=REG[0]<<0;
      10'h1d5: data = 32'h8c420000; // 00400754: LW, REG[2]<=RAM[REG[2]+0];
      10'h1d6: data = 32'h00000000; // 00400758: SLL, REG[0]<=REG[0]<<0;
      10'h1d7: data = 32'h2c420020; // 0040075c: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h1d8: data = 32'h14400010; // 00400760: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h1d9: data = 32'h00000000; // 00400764: SLL, REG[0]<=REG[0]<<0;
      10'h1da: data = 32'h8fc20008; // 00400768: LW, REG[2]<=RAM[REG[30]+8];
      10'h1db: data = 32'h00000000; // 0040076c: SLL, REG[0]<=REG[0]<<0;
      10'h1dc: data = 32'h8c420000; // 00400770: LW, REG[2]<=RAM[REG[2]+0];
      10'h1dd: data = 32'h00000000; // 00400774: SLL, REG[0]<=REG[0]<<0;
      10'h1de: data = 32'h2c420030; // 00400778: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h1df: data = 32'h10400009; // 0040077c: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h1e0: data = 32'h00000000; // 00400780: SLL, REG[0]<=REG[0]<<0;
      10'h1e1: data = 32'h8fc20008; // 00400784: LW, REG[2]<=RAM[REG[30]+8];
      10'h1e2: data = 32'h00000000; // 00400788: SLL, REG[0]<=REG[0]<<0;
      10'h1e3: data = 32'h8c430000; // 0040078c: LW, REG[3]<=RAM[REG[2]+0];
      10'h1e4: data = 32'h8fc20008; // 00400790: LW, REG[2]<=RAM[REG[30]+8];
      10'h1e5: data = 32'h00000000; // 00400794: SLL, REG[0]<=REG[0]<<0;
      10'h1e6: data = 32'hac430000; // 00400798: SW, RAM[REG[2]+0]<=REG[3];
      10'h1e7: data = 32'h08100223; // 0040079c: J, PC<=0x00100223*4(=0x0040088c);
      10'h1e8: data = 32'h00000000; // 004007a0: SLL, REG[0]<=REG[0]<<0;
      10'h1e9: data = 32'h8fc20008; // 004007a4: LW, REG[2]<=RAM[REG[30]+8];
      10'h1ea: data = 32'h00000000; // 004007a8: SLL, REG[0]<=REG[0]<<0;
      10'h1eb: data = 32'h8c430000; // 004007ac: LW, REG[3]<=RAM[REG[2]+0];
      10'h1ec: data = 32'h2402003a; // 004007b0: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h1ed: data = 32'h14620006; // 004007b4: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1ee: data = 32'h00000000; // 004007b8: SLL, REG[0]<=REG[0]<<0;
      10'h1ef: data = 32'h8fc30008; // 004007bc: LW, REG[3]<=RAM[REG[30]+8];
      10'h1f0: data = 32'h2402003f; // 004007c0: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h1f1: data = 32'hac620000; // 004007c4: SW, RAM[REG[3]+0]<=REG[2];
      10'h1f2: data = 32'h08100223; // 004007c8: J, PC<=0x00100223*4(=0x0040088c);
      10'h1f3: data = 32'h00000000; // 004007cc: SLL, REG[0]<=REG[0]<<0;
      10'h1f4: data = 32'h8fc20008; // 004007d0: LW, REG[2]<=RAM[REG[30]+8];
      10'h1f5: data = 32'h00000000; // 004007d4: SLL, REG[0]<=REG[0]<<0;
      10'h1f6: data = 32'h8c430000; // 004007d8: LW, REG[3]<=RAM[REG[2]+0];
      10'h1f7: data = 32'h2402003b; // 004007dc: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h1f8: data = 32'h14620006; // 004007e0: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1f9: data = 32'h00000000; // 004007e4: SLL, REG[0]<=REG[0]<<0;
      10'h1fa: data = 32'h8fc30008; // 004007e8: LW, REG[3]<=RAM[REG[30]+8];
      10'h1fb: data = 32'h2402003d; // 004007ec: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h1fc: data = 32'hac620000; // 004007f0: SW, RAM[REG[3]+0]<=REG[2];
      10'h1fd: data = 32'h08100223; // 004007f4: J, PC<=0x00100223*4(=0x0040088c);
      10'h1fe: data = 32'h00000000; // 004007f8: SLL, REG[0]<=REG[0]<<0;
      10'h1ff: data = 32'h8fc20008; // 004007fc: LW, REG[2]<=RAM[REG[30]+8];
      10'h200: data = 32'h00000000; // 00400800: SLL, REG[0]<=REG[0]<<0;
      10'h201: data = 32'h8c430000; // 00400804: LW, REG[3]<=RAM[REG[2]+0];
      10'h202: data = 32'h2402003c; // 00400808: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h203: data = 32'h14620006; // 0040080c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h204: data = 32'h00000000; // 00400810: SLL, REG[0]<=REG[0]<<0;
      10'h205: data = 32'h8fc30008; // 00400814: LW, REG[3]<=RAM[REG[30]+8];
      10'h206: data = 32'h2402003b; // 00400818: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h207: data = 32'hac620000; // 0040081c: SW, RAM[REG[3]+0]<=REG[2];
      10'h208: data = 32'h08100223; // 00400820: J, PC<=0x00100223*4(=0x0040088c);
      10'h209: data = 32'h00000000; // 00400824: SLL, REG[0]<=REG[0]<<0;
      10'h20a: data = 32'h8fc20008; // 00400828: LW, REG[2]<=RAM[REG[30]+8];
      10'h20b: data = 32'h00000000; // 0040082c: SLL, REG[0]<=REG[0]<<0;
      10'h20c: data = 32'h8c430000; // 00400830: LW, REG[3]<=RAM[REG[2]+0];
      10'h20d: data = 32'h2402003d; // 00400834: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h20e: data = 32'h14620006; // 00400838: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h20f: data = 32'h00000000; // 0040083c: SLL, REG[0]<=REG[0]<<0;
      10'h210: data = 32'h8fc30008; // 00400840: LW, REG[3]<=RAM[REG[30]+8];
      10'h211: data = 32'h2402003a; // 00400844: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h212: data = 32'hac620000; // 00400848: SW, RAM[REG[3]+0]<=REG[2];
      10'h213: data = 32'h08100223; // 0040084c: J, PC<=0x00100223*4(=0x0040088c);
      10'h214: data = 32'h00000000; // 00400850: SLL, REG[0]<=REG[0]<<0;
      10'h215: data = 32'h8fc20008; // 00400854: LW, REG[2]<=RAM[REG[30]+8];
      10'h216: data = 32'h00000000; // 00400858: SLL, REG[0]<=REG[0]<<0;
      10'h217: data = 32'h8c430000; // 0040085c: LW, REG[3]<=RAM[REG[2]+0];
      10'h218: data = 32'h2402003e; // 00400860: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h219: data = 32'h14620006; // 00400864: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h21a: data = 32'h00000000; // 00400868: SLL, REG[0]<=REG[0]<<0;
      10'h21b: data = 32'h8fc30008; // 0040086c: LW, REG[3]<=RAM[REG[30]+8];
      10'h21c: data = 32'h2402000a; // 00400870: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h21d: data = 32'hac620000; // 00400874: SW, RAM[REG[3]+0]<=REG[2];
      10'h21e: data = 32'h08100223; // 00400878: J, PC<=0x00100223*4(=0x0040088c);
      10'h21f: data = 32'h00000000; // 0040087c: SLL, REG[0]<=REG[0]<<0;
      10'h220: data = 32'h8fc30008; // 00400880: LW, REG[3]<=RAM[REG[30]+8];
      10'h221: data = 32'h24020040; // 00400884: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h222: data = 32'hac620000; // 00400888: SW, RAM[REG[3]+0]<=REG[2];
      10'h223: data = 32'h24020308; // 0040088c: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h224: data = 32'hac400000; // 00400890: SW, RAM[REG[2]+0]<=REG[0];
      10'h225: data = 32'h24030308; // 00400894: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h226: data = 32'h24020001; // 00400898: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h227: data = 32'hac620000; // 0040089c: SW, RAM[REG[3]+0]<=REG[2];
      10'h228: data = 32'h8fc20008; // 004008a0: LW, REG[2]<=RAM[REG[30]+8];
      10'h229: data = 32'h00000000; // 004008a4: SLL, REG[0]<=REG[0]<<0;
      10'h22a: data = 32'h24420004; // 004008a8: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h22b: data = 32'hafc20008; // 004008ac: SW, RAM[REG[30]+8]<=REG[2];
      10'h22c: data = 32'h24020310; // 004008b0: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h22d: data = 32'h8c430000; // 004008b4: LW, REG[3]<=RAM[REG[2]+0];
      10'h22e: data = 32'h8fc20008; // 004008b8: LW, REG[2]<=RAM[REG[30]+8];
      10'h22f: data = 32'h00000000; // 004008bc: SLL, REG[0]<=REG[0]<<0;
      10'h230: data = 32'hac430000; // 004008c0: SW, RAM[REG[2]+0]<=REG[3];
      10'h231: data = 32'h8fc20008; // 004008c4: LW, REG[2]<=RAM[REG[30]+8];
      10'h232: data = 32'h00000000; // 004008c8: SLL, REG[0]<=REG[0]<<0;
      10'h233: data = 32'h8c430000; // 004008cc: LW, REG[3]<=RAM[REG[2]+0];
      10'h234: data = 32'h2402003e; // 004008d0: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h235: data = 32'h1462ff4f; // 004008d4: BNE, PC<=(REG[3] != REG[2])?PC+4+65359*4:PC+4;
      10'h236: data = 32'h00000000; // 004008d8: SLL, REG[0]<=REG[0]<<0;
      10'h237: data = 32'h8fc20008; // 004008dc: LW, REG[2]<=RAM[REG[30]+8];
      10'h238: data = 32'h00000000; // 004008e0: SLL, REG[0]<=REG[0]<<0;
      10'h239: data = 32'hac400000; // 004008e4: SW, RAM[REG[2]+0]<=REG[0];
      10'h23a: data = 32'h24020308; // 004008e8: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h23b: data = 32'hac400000; // 004008ec: SW, RAM[REG[2]+0]<=REG[0];
      10'h23c: data = 32'h2402030c; // 004008f0: ADDIU, REG[2]<=REG[0]+780(=0x0000030c);
      10'h23d: data = 32'hac400000; // 004008f4: SW, RAM[REG[2]+0]<=REG[0];
      10'h23e: data = 32'h24030308; // 004008f8: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h23f: data = 32'h24020001; // 004008fc: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h240: data = 32'hac620000; // 00400900: SW, RAM[REG[3]+0]<=REG[2];
      10'h241: data = 32'h24020308; // 00400904: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h242: data = 32'hac400000; // 00400908: SW, RAM[REG[2]+0]<=REG[0];
      10'h243: data = 32'h03c0e821; // 0040090c: ADDU, REG[29]<=REG[30]+REG[0];
      10'h244: data = 32'h8fbe0000; // 00400910: LW, REG[30]<=RAM[REG[29]+0];
      10'h245: data = 32'h27bd0008; // 00400914: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h246: data = 32'h03e00008; // 00400918: JR, PC<=REG[31];
      10'h247: data = 32'h00000000; // 0040091c: SLL, REG[0]<=REG[0]<<0;
      10'h248: data = 32'h27bdfff8; // 00400920: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h249: data = 32'hafbe0000; // 00400924: SW, RAM[REG[29]+0]<=REG[30];
      10'h24a: data = 32'h03a0f021; // 00400928: ADDU, REG[30]<=REG[29]+REG[0];
      10'h24b: data = 32'hafc40008; // 0040092c: SW, RAM[REG[30]+8]<=REG[4];
      10'h24c: data = 32'h0810030a; // 00400930: J, PC<=0x0010030a*4(=0x00400c28);
      10'h24d: data = 32'h00000000; // 00400934: SLL, REG[0]<=REG[0]<<0;
      10'h24e: data = 32'h24020300; // 00400938: ADDIU, REG[2]<=REG[0]+768(=0x00000300);
      10'h24f: data = 32'hac400000; // 0040093c: SW, RAM[REG[2]+0]<=REG[0];
      10'h250: data = 32'h8fc20008; // 00400940: LW, REG[2]<=RAM[REG[30]+8];
      10'h251: data = 32'h00000000; // 00400944: SLL, REG[0]<=REG[0]<<0;
      10'h252: data = 32'h8c420000; // 00400948: LW, REG[2]<=RAM[REG[2]+0];
      10'h253: data = 32'h00000000; // 0040094c: SLL, REG[0]<=REG[0]<<0;
      10'h254: data = 32'h2c420041; // 00400950: SLTIU, REG[2]<=(REG[2]<65(=0x00000041))?1:0;
      10'h255: data = 32'h14400011; // 00400954: BNE, PC<=(REG[2] != REG[0])?PC+4+17*4:PC+4;
      10'h256: data = 32'h00000000; // 00400958: SLL, REG[0]<=REG[0]<<0;
      10'h257: data = 32'h8fc20008; // 0040095c: LW, REG[2]<=RAM[REG[30]+8];
      10'h258: data = 32'h00000000; // 00400960: SLL, REG[0]<=REG[0]<<0;
      10'h259: data = 32'h8c420000; // 00400964: LW, REG[2]<=RAM[REG[2]+0];
      10'h25a: data = 32'h00000000; // 00400968: SLL, REG[0]<=REG[0]<<0;
      10'h25b: data = 32'h2c42005b; // 0040096c: SLTIU, REG[2]<=(REG[2]<91(=0x0000005b))?1:0;
      10'h25c: data = 32'h1040000a; // 00400970: BEQ, PC<=(REG[2] == REG[0])?PC+4+10*4:PC+4;
      10'h25d: data = 32'h00000000; // 00400974: SLL, REG[0]<=REG[0]<<0;
      10'h25e: data = 32'h24030304; // 00400978: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h25f: data = 32'h8fc20008; // 0040097c: LW, REG[2]<=RAM[REG[30]+8];
      10'h260: data = 32'h00000000; // 00400980: SLL, REG[0]<=REG[0]<<0;
      10'h261: data = 32'h8c420000; // 00400984: LW, REG[2]<=RAM[REG[2]+0];
      10'h262: data = 32'h00000000; // 00400988: SLL, REG[0]<=REG[0]<<0;
      10'h263: data = 32'h2442ffc0; // 0040098c: ADDIU, REG[2]<=REG[2]+65472(=0x0000ffc0);
      10'h264: data = 32'hac620000; // 00400990: SW, RAM[REG[3]+0]<=REG[2];
      10'h265: data = 32'h08100303; // 00400994: J, PC<=0x00100303*4(=0x00400c0c);
      10'h266: data = 32'h00000000; // 00400998: SLL, REG[0]<=REG[0]<<0;
      10'h267: data = 32'h8fc20008; // 0040099c: LW, REG[2]<=RAM[REG[30]+8];
      10'h268: data = 32'h00000000; // 004009a0: SLL, REG[0]<=REG[0]<<0;
      10'h269: data = 32'h8c420000; // 004009a4: LW, REG[2]<=RAM[REG[2]+0];
      10'h26a: data = 32'h00000000; // 004009a8: SLL, REG[0]<=REG[0]<<0;
      10'h26b: data = 32'h2c420061; // 004009ac: SLTIU, REG[2]<=(REG[2]<97(=0x00000061))?1:0;
      10'h26c: data = 32'h14400011; // 004009b0: BNE, PC<=(REG[2] != REG[0])?PC+4+17*4:PC+4;
      10'h26d: data = 32'h00000000; // 004009b4: SLL, REG[0]<=REG[0]<<0;
      10'h26e: data = 32'h8fc20008; // 004009b8: LW, REG[2]<=RAM[REG[30]+8];
      10'h26f: data = 32'h00000000; // 004009bc: SLL, REG[0]<=REG[0]<<0;
      10'h270: data = 32'h8c420000; // 004009c0: LW, REG[2]<=RAM[REG[2]+0];
      10'h271: data = 32'h00000000; // 004009c4: SLL, REG[0]<=REG[0]<<0;
      10'h272: data = 32'h2c42007b; // 004009c8: SLTIU, REG[2]<=(REG[2]<123(=0x0000007b))?1:0;
      10'h273: data = 32'h1040000a; // 004009cc: BEQ, PC<=(REG[2] == REG[0])?PC+4+10*4:PC+4;
      10'h274: data = 32'h00000000; // 004009d0: SLL, REG[0]<=REG[0]<<0;
      10'h275: data = 32'h24030304; // 004009d4: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h276: data = 32'h8fc20008; // 004009d8: LW, REG[2]<=RAM[REG[30]+8];
      10'h277: data = 32'h00000000; // 004009dc: SLL, REG[0]<=REG[0]<<0;
      10'h278: data = 32'h8c420000; // 004009e0: LW, REG[2]<=RAM[REG[2]+0];
      10'h279: data = 32'h00000000; // 004009e4: SLL, REG[0]<=REG[0]<<0;
      10'h27a: data = 32'h2442ffa0; // 004009e8: ADDIU, REG[2]<=REG[2]+65440(=0x0000ffa0);
      10'h27b: data = 32'hac620000; // 004009ec: SW, RAM[REG[3]+0]<=REG[2];
      10'h27c: data = 32'h08100303; // 004009f0: J, PC<=0x00100303*4(=0x00400c0c);
      10'h27d: data = 32'h00000000; // 004009f4: SLL, REG[0]<=REG[0]<<0;
      10'h27e: data = 32'h8fc20008; // 004009f8: LW, REG[2]<=RAM[REG[30]+8];
      10'h27f: data = 32'h00000000; // 004009fc: SLL, REG[0]<=REG[0]<<0;
      10'h280: data = 32'h8c420000; // 00400a00: LW, REG[2]<=RAM[REG[2]+0];
      10'h281: data = 32'h00000000; // 00400a04: SLL, REG[0]<=REG[0]<<0;
      10'h282: data = 32'h2c420030; // 00400a08: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h283: data = 32'h14400010; // 00400a0c: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h284: data = 32'h00000000; // 00400a10: SLL, REG[0]<=REG[0]<<0;
      10'h285: data = 32'h8fc20008; // 00400a14: LW, REG[2]<=RAM[REG[30]+8];
      10'h286: data = 32'h00000000; // 00400a18: SLL, REG[0]<=REG[0]<<0;
      10'h287: data = 32'h8c420000; // 00400a1c: LW, REG[2]<=RAM[REG[2]+0];
      10'h288: data = 32'h00000000; // 00400a20: SLL, REG[0]<=REG[0]<<0;
      10'h289: data = 32'h2c42003a; // 00400a24: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h28a: data = 32'h10400009; // 00400a28: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h28b: data = 32'h00000000; // 00400a2c: SLL, REG[0]<=REG[0]<<0;
      10'h28c: data = 32'h24020304; // 00400a30: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h28d: data = 32'h8fc30008; // 00400a34: LW, REG[3]<=RAM[REG[30]+8];
      10'h28e: data = 32'h00000000; // 00400a38: SLL, REG[0]<=REG[0]<<0;
      10'h28f: data = 32'h8c630000; // 00400a3c: LW, REG[3]<=RAM[REG[3]+0];
      10'h290: data = 32'h00000000; // 00400a40: SLL, REG[0]<=REG[0]<<0;
      10'h291: data = 32'hac430000; // 00400a44: SW, RAM[REG[2]+0]<=REG[3];
      10'h292: data = 32'h08100303; // 00400a48: J, PC<=0x00100303*4(=0x00400c0c);
      10'h293: data = 32'h00000000; // 00400a4c: SLL, REG[0]<=REG[0]<<0;
      10'h294: data = 32'h8fc20008; // 00400a50: LW, REG[2]<=RAM[REG[30]+8];
      10'h295: data = 32'h00000000; // 00400a54: SLL, REG[0]<=REG[0]<<0;
      10'h296: data = 32'h8c430000; // 00400a58: LW, REG[3]<=RAM[REG[2]+0];
      10'h297: data = 32'h24020040; // 00400a5c: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h298: data = 32'h14620005; // 00400a60: BNE, PC<=(REG[3] != REG[2])?PC+4+5*4:PC+4;
      10'h299: data = 32'h00000000; // 00400a64: SLL, REG[0]<=REG[0]<<0;
      10'h29a: data = 32'h24020304; // 00400a68: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h29b: data = 32'hac400000; // 00400a6c: SW, RAM[REG[2]+0]<=REG[0];
      10'h29c: data = 32'h08100303; // 00400a70: J, PC<=0x00100303*4(=0x00400c0c);
      10'h29d: data = 32'h00000000; // 00400a74: SLL, REG[0]<=REG[0]<<0;
      10'h29e: data = 32'h8fc20008; // 00400a78: LW, REG[2]<=RAM[REG[30]+8];
      10'h29f: data = 32'h00000000; // 00400a7c: SLL, REG[0]<=REG[0]<<0;
      10'h2a0: data = 32'h8c430000; // 00400a80: LW, REG[3]<=RAM[REG[2]+0];
      10'h2a1: data = 32'h2402005b; // 00400a84: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h2a2: data = 32'h14620006; // 00400a88: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2a3: data = 32'h00000000; // 00400a8c: SLL, REG[0]<=REG[0]<<0;
      10'h2a4: data = 32'h24030304; // 00400a90: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h2a5: data = 32'h2402001b; // 00400a94: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h2a6: data = 32'hac620000; // 00400a98: SW, RAM[REG[3]+0]<=REG[2];
      10'h2a7: data = 32'h08100303; // 00400a9c: J, PC<=0x00100303*4(=0x00400c0c);
      10'h2a8: data = 32'h00000000; // 00400aa0: SLL, REG[0]<=REG[0]<<0;
      10'h2a9: data = 32'h8fc20008; // 00400aa4: LW, REG[2]<=RAM[REG[30]+8];
      10'h2aa: data = 32'h00000000; // 00400aa8: SLL, REG[0]<=REG[0]<<0;
      10'h2ab: data = 32'h8c430000; // 00400aac: LW, REG[3]<=RAM[REG[2]+0];
      10'h2ac: data = 32'h2402005d; // 00400ab0: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h2ad: data = 32'h14620006; // 00400ab4: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2ae: data = 32'h00000000; // 00400ab8: SLL, REG[0]<=REG[0]<<0;
      10'h2af: data = 32'h24030304; // 00400abc: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h2b0: data = 32'h2402001d; // 00400ac0: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h2b1: data = 32'hac620000; // 00400ac4: SW, RAM[REG[3]+0]<=REG[2];
      10'h2b2: data = 32'h08100303; // 00400ac8: J, PC<=0x00100303*4(=0x00400c0c);
      10'h2b3: data = 32'h00000000; // 00400acc: SLL, REG[0]<=REG[0]<<0;
      10'h2b4: data = 32'h8fc20008; // 00400ad0: LW, REG[2]<=RAM[REG[30]+8];
      10'h2b5: data = 32'h00000000; // 00400ad4: SLL, REG[0]<=REG[0]<<0;
      10'h2b6: data = 32'h8c420000; // 00400ad8: LW, REG[2]<=RAM[REG[2]+0];
      10'h2b7: data = 32'h00000000; // 00400adc: SLL, REG[0]<=REG[0]<<0;
      10'h2b8: data = 32'h2c420020; // 00400ae0: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h2b9: data = 32'h14400010; // 00400ae4: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h2ba: data = 32'h00000000; // 00400ae8: SLL, REG[0]<=REG[0]<<0;
      10'h2bb: data = 32'h8fc20008; // 00400aec: LW, REG[2]<=RAM[REG[30]+8];
      10'h2bc: data = 32'h00000000; // 00400af0: SLL, REG[0]<=REG[0]<<0;
      10'h2bd: data = 32'h8c420000; // 00400af4: LW, REG[2]<=RAM[REG[2]+0];
      10'h2be: data = 32'h00000000; // 00400af8: SLL, REG[0]<=REG[0]<<0;
      10'h2bf: data = 32'h2c420030; // 00400afc: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h2c0: data = 32'h10400009; // 00400b00: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h2c1: data = 32'h00000000; // 00400b04: SLL, REG[0]<=REG[0]<<0;
      10'h2c2: data = 32'h24020304; // 00400b08: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h2c3: data = 32'h8fc30008; // 00400b0c: LW, REG[3]<=RAM[REG[30]+8];
      10'h2c4: data = 32'h00000000; // 00400b10: SLL, REG[0]<=REG[0]<<0;
      10'h2c5: data = 32'h8c630000; // 00400b14: LW, REG[3]<=RAM[REG[3]+0];
      10'h2c6: data = 32'h00000000; // 00400b18: SLL, REG[0]<=REG[0]<<0;
      10'h2c7: data = 32'hac430000; // 00400b1c: SW, RAM[REG[2]+0]<=REG[3];
      10'h2c8: data = 32'h08100303; // 00400b20: J, PC<=0x00100303*4(=0x00400c0c);
      10'h2c9: data = 32'h00000000; // 00400b24: SLL, REG[0]<=REG[0]<<0;
      10'h2ca: data = 32'h8fc20008; // 00400b28: LW, REG[2]<=RAM[REG[30]+8];
      10'h2cb: data = 32'h00000000; // 00400b2c: SLL, REG[0]<=REG[0]<<0;
      10'h2cc: data = 32'h8c430000; // 00400b30: LW, REG[3]<=RAM[REG[2]+0];
      10'h2cd: data = 32'h2402003f; // 00400b34: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h2ce: data = 32'h14620006; // 00400b38: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2cf: data = 32'h00000000; // 00400b3c: SLL, REG[0]<=REG[0]<<0;
      10'h2d0: data = 32'h24030304; // 00400b40: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h2d1: data = 32'h2402003a; // 00400b44: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h2d2: data = 32'hac620000; // 00400b48: SW, RAM[REG[3]+0]<=REG[2];
      10'h2d3: data = 32'h08100303; // 00400b4c: J, PC<=0x00100303*4(=0x00400c0c);
      10'h2d4: data = 32'h00000000; // 00400b50: SLL, REG[0]<=REG[0]<<0;
      10'h2d5: data = 32'h8fc20008; // 00400b54: LW, REG[2]<=RAM[REG[30]+8];
      10'h2d6: data = 32'h00000000; // 00400b58: SLL, REG[0]<=REG[0]<<0;
      10'h2d7: data = 32'h8c430000; // 00400b5c: LW, REG[3]<=RAM[REG[2]+0];
      10'h2d8: data = 32'h2402003d; // 00400b60: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h2d9: data = 32'h14620006; // 00400b64: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2da: data = 32'h00000000; // 00400b68: SLL, REG[0]<=REG[0]<<0;
      10'h2db: data = 32'h24030304; // 00400b6c: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h2dc: data = 32'h2402003b; // 00400b70: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h2dd: data = 32'hac620000; // 00400b74: SW, RAM[REG[3]+0]<=REG[2];
      10'h2de: data = 32'h08100303; // 00400b78: J, PC<=0x00100303*4(=0x00400c0c);
      10'h2df: data = 32'h00000000; // 00400b7c: SLL, REG[0]<=REG[0]<<0;
      10'h2e0: data = 32'h8fc20008; // 00400b80: LW, REG[2]<=RAM[REG[30]+8];
      10'h2e1: data = 32'h00000000; // 00400b84: SLL, REG[0]<=REG[0]<<0;
      10'h2e2: data = 32'h8c430000; // 00400b88: LW, REG[3]<=RAM[REG[2]+0];
      10'h2e3: data = 32'h2402003b; // 00400b8c: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h2e4: data = 32'h14620006; // 00400b90: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2e5: data = 32'h00000000; // 00400b94: SLL, REG[0]<=REG[0]<<0;
      10'h2e6: data = 32'h24030304; // 00400b98: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h2e7: data = 32'h2402003c; // 00400b9c: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h2e8: data = 32'hac620000; // 00400ba0: SW, RAM[REG[3]+0]<=REG[2];
      10'h2e9: data = 32'h08100303; // 00400ba4: J, PC<=0x00100303*4(=0x00400c0c);
      10'h2ea: data = 32'h00000000; // 00400ba8: SLL, REG[0]<=REG[0]<<0;
      10'h2eb: data = 32'h8fc20008; // 00400bac: LW, REG[2]<=RAM[REG[30]+8];
      10'h2ec: data = 32'h00000000; // 00400bb0: SLL, REG[0]<=REG[0]<<0;
      10'h2ed: data = 32'h8c430000; // 00400bb4: LW, REG[3]<=RAM[REG[2]+0];
      10'h2ee: data = 32'h2402003a; // 00400bb8: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h2ef: data = 32'h14620006; // 00400bbc: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2f0: data = 32'h00000000; // 00400bc0: SLL, REG[0]<=REG[0]<<0;
      10'h2f1: data = 32'h24030304; // 00400bc4: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h2f2: data = 32'h2402003d; // 00400bc8: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h2f3: data = 32'hac620000; // 00400bcc: SW, RAM[REG[3]+0]<=REG[2];
      10'h2f4: data = 32'h08100303; // 00400bd0: J, PC<=0x00100303*4(=0x00400c0c);
      10'h2f5: data = 32'h00000000; // 00400bd4: SLL, REG[0]<=REG[0]<<0;
      10'h2f6: data = 32'h8fc20008; // 00400bd8: LW, REG[2]<=RAM[REG[30]+8];
      10'h2f7: data = 32'h00000000; // 00400bdc: SLL, REG[0]<=REG[0]<<0;
      10'h2f8: data = 32'h8c430000; // 00400be0: LW, REG[3]<=RAM[REG[2]+0];
      10'h2f9: data = 32'h2402000a; // 00400be4: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h2fa: data = 32'h14620006; // 00400be8: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2fb: data = 32'h00000000; // 00400bec: SLL, REG[0]<=REG[0]<<0;
      10'h2fc: data = 32'h24030304; // 00400bf0: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h2fd: data = 32'h2402003e; // 00400bf4: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h2fe: data = 32'hac620000; // 00400bf8: SW, RAM[REG[3]+0]<=REG[2];
      10'h2ff: data = 32'h08100303; // 00400bfc: J, PC<=0x00100303*4(=0x00400c0c);
      10'h300: data = 32'h00000000; // 00400c00: SLL, REG[0]<=REG[0]<<0;
      10'h301: data = 32'h24020304; // 00400c04: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h302: data = 32'hac400000; // 00400c08: SW, RAM[REG[2]+0]<=REG[0];
      10'h303: data = 32'h24030300; // 00400c0c: ADDIU, REG[3]<=REG[0]+768(=0x00000300);
      10'h304: data = 32'h24020001; // 00400c10: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h305: data = 32'hac620000; // 00400c14: SW, RAM[REG[3]+0]<=REG[2];
      10'h306: data = 32'h8fc20008; // 00400c18: LW, REG[2]<=RAM[REG[30]+8];
      10'h307: data = 32'h00000000; // 00400c1c: SLL, REG[0]<=REG[0]<<0;
      10'h308: data = 32'h24420004; // 00400c20: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h309: data = 32'hafc20008; // 00400c24: SW, RAM[REG[30]+8]<=REG[2];
      10'h30a: data = 32'h8fc20008; // 00400c28: LW, REG[2]<=RAM[REG[30]+8];
      10'h30b: data = 32'h00000000; // 00400c2c: SLL, REG[0]<=REG[0]<<0;
      10'h30c: data = 32'h8c420000; // 00400c30: LW, REG[2]<=RAM[REG[2]+0];
      10'h30d: data = 32'h00000000; // 00400c34: SLL, REG[0]<=REG[0]<<0;
      10'h30e: data = 32'h1440ff3f; // 00400c38: BNE, PC<=(REG[2] != REG[0])?PC+4+65343*4:PC+4;
      10'h30f: data = 32'h00000000; // 00400c3c: SLL, REG[0]<=REG[0]<<0;
      10'h310: data = 32'h03c0e821; // 00400c40: ADDU, REG[29]<=REG[30]+REG[0];
      10'h311: data = 32'h8fbe0000; // 00400c44: LW, REG[30]<=RAM[REG[29]+0];
      10'h312: data = 32'h27bd0008; // 00400c48: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h313: data = 32'h03e00008; // 00400c4c: JR, PC<=REG[31];
      10'h314: data = 32'h00000000; // 00400c50: SLL, REG[0]<=REG[0]<<0;
      10'h315: data = 32'h00000000; // 00400c54: SLL, REG[0]<=REG[0]<<0;
      10'h316: data = 32'h00000000; // 00400c58: SLL, REG[0]<=REG[0]<<0;
      10'h317: data = 32'h00000000; // 00400c5c: SLL, REG[0]<=REG[0]<<0;
    endcase
  end

  assign rom_data = data;
endmodule
