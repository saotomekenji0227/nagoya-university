library verilog;
use verilog.vl_types.all;
entity test_mux21 is
end test_mux21;
