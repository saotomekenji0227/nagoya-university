/*                                 *
 * test_bcd1.v                     *
 * 1���BCD�����󥿤Υƥ��ȥ٥��      *
 *                                 */
 
`timescale 1ns / 1ns    // ���ߥ�졼������ñ�̻��� / ����
                                                // 1ns = 1/1000000000 sec
`include "bcd1.v"   // bcd1.v ���ɤ߹���
 
module test ;
  /*** bcd1 �������ͳ�Ǽ�ѤΥ쥸���� ****/
  reg reset, clk, x;

  /*** bcd1 �ν��ϴ�¬�Ѥο����� ****/
  wire [3:0] bcd1_out;

  /*** bcd1 �μ��β� ***/
   bcd1 bcd1a(clk, reset, x, bcd1_out);
 
  always begin
    #5      clk = ~clk;
  end
 
  always begin
    #15     x = ~x;
  end
 
  initial begin
    reset = 1; clk = 0; x = 0;

    // 20 ñ�̻���(20 ns)��
    #20 reset = 0;

    // ���� 20 ñ�̻���(20 ns)��
    #20 reset = 1;

    // ���� 1000 ñ�̻���(1000 ns)��, ��λ
    #1000 $finish;
  end
 
endmodule // test
