/*******************/
/* rom8x1024_sim.v */
/*******************/

//                  +----+
//  rom_addr[11:0]->|    |->rom_data[31:0]
//                  +----+

//
// ROM�ε��ҡ��������ߥ�졼������ѡ�
//

module rom8x1024_sim (rom_addr, rom_data);

  input   [11:0]  rom_addr;  // 12-bit ���ɥ쥹���ϥݡ���
  output  [31:0]  rom_data;  // 32-bit �ǡ������ϥݡ���

  reg     [31:0]  data;

  // Wire
  wire     [9:0]  word_addr; // 10-bit address, word

  assign word_addr = rom_addr[9:2];
   
  always @(word_addr) begin
    case (word_addr)
      10'h000: data = 32'he000001c; // 00400000: other type! opcode=56(10)
      10'h001: data = 32'h00000000; // 00400004: SLL, REG[0]<=REG[0]<<0;
      10'h002: data = 32'h00000000; // 00400008: SLL, REG[0]<=REG[0]<<0;
      10'h003: data = 32'h00000000; // 0040000c: SLL, REG[0]<=REG[0]<<0;
      10'h004: data = 32'h00000000; // 00400010: SLL, REG[0]<=REG[0]<<0;
      10'h005: data = 32'h004088b0; // 00400014: R type, unknown. func=48(10)
      10'h006: data = 32'h00000000; // 00400018: SLL, REG[0]<=REG[0]<<0;
      10'h007: data = 32'h00000000; // 0040001c: SLL, REG[0]<=REG[0]<<0;
      10'h008: data = 32'h27bdff98; // 00400020: ADDIU, REG[29]<=REG[29]+65432(=0x0000ff98);
      10'h009: data = 32'hafbf0064; // 00400024: SW, RAM[REG[29]+100]<=REG[31];
      10'h00a: data = 32'hafbe0060; // 00400028: SW, RAM[REG[29]+96]<=REG[30];
      10'h00b: data = 32'h03a0f021; // 0040002c: ADDU, REG[30]<=REG[29]+REG[0];
      10'h00c: data = 32'hafc00018; // 00400030: SW, RAM[REG[30]+24]<=REG[0];
      10'h00d: data = 32'h27c2001c; // 00400034: ADDIU, REG[2]<=REG[30]+28(=0x0000001c);
      10'h00e: data = 32'h00402021; // 00400038: ADDU, REG[4]<=REG[2]+REG[0];
      10'h00f: data = 32'h0c1000b9; // 0040003c: JAL, PC<=0x001000b9*4(=0x004002e4); REG[31]<=PC+4
      10'h010: data = 32'h00000000; // 00400040: SLL, REG[0]<=REG[0]<<0;
      10'h011: data = 32'h8fc3001c; // 00400044: LW, REG[3]<=RAM[REG[30]+28];
      10'h012: data = 32'h24020052; // 00400048: ADDIU, REG[2]<=REG[0]+82(=0x00000052);
      10'h013: data = 32'h14620004; // 0040004c: BNE, PC<=(REG[3] != REG[2])?PC+4+4*4:PC+4;
      10'h014: data = 32'h00000000; // 00400050: SLL, REG[0]<=REG[0]<<0;
      10'h015: data = 32'hafc00018; // 00400054: SW, RAM[REG[30]+24]<=REG[0];
      10'h016: data = 32'h08100026; // 00400058: J, PC<=0x00100026*4(=0x00400098);
      10'h017: data = 32'h00000000; // 0040005c: SLL, REG[0]<=REG[0]<<0;
      10'h018: data = 32'h8fc3001c; // 00400060: LW, REG[3]<=RAM[REG[30]+28];
      10'h019: data = 32'h2402004c; // 00400064: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h01a: data = 32'h14620005; // 00400068: BNE, PC<=(REG[3] != REG[2])?PC+4+5*4:PC+4;
      10'h01b: data = 32'h00000000; // 0040006c: SLL, REG[0]<=REG[0]<<0;
      10'h01c: data = 32'h24020001; // 00400070: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h01d: data = 32'hafc20018; // 00400074: SW, RAM[REG[30]+24]<=REG[2];
      10'h01e: data = 32'h08100026; // 00400078: J, PC<=0x00100026*4(=0x00400098);
      10'h01f: data = 32'h00000000; // 0040007c: SLL, REG[0]<=REG[0]<<0;
      10'h020: data = 32'h8fc3001c; // 00400080: LW, REG[3]<=RAM[REG[30]+28];
      10'h021: data = 32'h24020053; // 00400084: ADDIU, REG[2]<=REG[0]+83(=0x00000053);
      10'h022: data = 32'h14620003; // 00400088: BNE, PC<=(REG[3] != REG[2])?PC+4+3*4:PC+4;
      10'h023: data = 32'h00000000; // 0040008c: SLL, REG[0]<=REG[0]<<0;
      10'h024: data = 32'h24020002; // 00400090: ADDIU, REG[2]<=REG[0]+2(=0x00000002);
      10'h025: data = 32'hafc20018; // 00400094: SW, RAM[REG[30]+24]<=REG[2];
      10'h026: data = 32'h27c2001c; // 00400098: ADDIU, REG[2]<=REG[30]+28(=0x0000001c);
      10'h027: data = 32'h00402021; // 0040009c: ADDU, REG[4]<=REG[2]+REG[0];
      10'h028: data = 32'h0c1000b9; // 004000a0: JAL, PC<=0x001000b9*4(=0x004002e4); REG[31]<=PC+4
      10'h029: data = 32'h00000000; // 004000a4: SLL, REG[0]<=REG[0]<<0;
      10'h02a: data = 32'h27c2001c; // 004000a8: ADDIU, REG[2]<=REG[30]+28(=0x0000001c);
      10'h02b: data = 32'h00402021; // 004000ac: ADDU, REG[4]<=REG[2]+REG[0];
      10'h02c: data = 32'h0c10019b; // 004000b0: JAL, PC<=0x0010019b*4(=0x0040066c); REG[31]<=PC+4
      10'h02d: data = 32'h00000000; // 004000b4: SLL, REG[0]<=REG[0]<<0;
      10'h02e: data = 32'hafc20010; // 004000b8: SW, RAM[REG[30]+16]<=REG[2];
      10'h02f: data = 32'h8fc20018; // 004000bc: LW, REG[2]<=RAM[REG[30]+24];
      10'h030: data = 32'h00000000; // 004000c0: SLL, REG[0]<=REG[0]<<0;
      10'h031: data = 32'h14400012; // 004000c4: BNE, PC<=(REG[2] != REG[0])?PC+4+18*4:PC+4;
      10'h032: data = 32'h00000000; // 004000c8: SLL, REG[0]<=REG[0]<<0;
      10'h033: data = 32'hafc00014; // 004000cc: SW, RAM[REG[30]+20]<=REG[0];
      10'h034: data = 32'h0810003c; // 004000d0: J, PC<=0x0010003c*4(=0x004000f0);
      10'h035: data = 32'h00000000; // 004000d4: SLL, REG[0]<=REG[0]<<0;
      10'h036: data = 32'h0c10006a; // 004000d8: JAL, PC<=0x0010006a*4(=0x004001a8); REG[31]<=PC+4
      10'h037: data = 32'h00000000; // 004000dc: SLL, REG[0]<=REG[0]<<0;
      10'h038: data = 32'h8fc20014; // 004000e0: LW, REG[2]<=RAM[REG[30]+20];
      10'h039: data = 32'h00000000; // 004000e4: SLL, REG[0]<=REG[0]<<0;
      10'h03a: data = 32'h24420001; // 004000e8: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h03b: data = 32'hafc20014; // 004000ec: SW, RAM[REG[30]+20]<=REG[2];
      10'h03c: data = 32'h8fc20014; // 004000f0: LW, REG[2]<=RAM[REG[30]+20];
      10'h03d: data = 32'h8fc30010; // 004000f4: LW, REG[3]<=RAM[REG[30]+16];
      10'h03e: data = 32'h00000000; // 004000f8: SLL, REG[0]<=REG[0]<<0;
      10'h03f: data = 32'h0043102b; // 004000fc: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h040: data = 32'h1440fff5; // 00400100: BNE, PC<=(REG[2] != REG[0])?PC+4+65525*4:PC+4;
      10'h041: data = 32'h00000000; // 00400104: SLL, REG[0]<=REG[0]<<0;
      10'h042: data = 32'h0810000d; // 00400108: J, PC<=0x0010000d*4(=0x00400034);
      10'h043: data = 32'h00000000; // 0040010c: SLL, REG[0]<=REG[0]<<0;
      10'h044: data = 32'h8fc30018; // 00400110: LW, REG[3]<=RAM[REG[30]+24];
      10'h045: data = 32'h24020001; // 00400114: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h046: data = 32'h14620012; // 00400118: BNE, PC<=(REG[3] != REG[2])?PC+4+18*4:PC+4;
      10'h047: data = 32'h00000000; // 0040011c: SLL, REG[0]<=REG[0]<<0;
      10'h048: data = 32'hafc00014; // 00400120: SW, RAM[REG[30]+20]<=REG[0];
      10'h049: data = 32'h08100051; // 00400124: J, PC<=0x00100051*4(=0x00400144);
      10'h04a: data = 32'h00000000; // 00400128: SLL, REG[0]<=REG[0]<<0;
      10'h04b: data = 32'h0c100080; // 0040012c: JAL, PC<=0x00100080*4(=0x00400200); REG[31]<=PC+4
      10'h04c: data = 32'h00000000; // 00400130: SLL, REG[0]<=REG[0]<<0;
      10'h04d: data = 32'h8fc20014; // 00400134: LW, REG[2]<=RAM[REG[30]+20];
      10'h04e: data = 32'h00000000; // 00400138: SLL, REG[0]<=REG[0]<<0;
      10'h04f: data = 32'h24420001; // 0040013c: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h050: data = 32'hafc20014; // 00400140: SW, RAM[REG[30]+20]<=REG[2];
      10'h051: data = 32'h8fc20014; // 00400144: LW, REG[2]<=RAM[REG[30]+20];
      10'h052: data = 32'h8fc30010; // 00400148: LW, REG[3]<=RAM[REG[30]+16];
      10'h053: data = 32'h00000000; // 0040014c: SLL, REG[0]<=REG[0]<<0;
      10'h054: data = 32'h0043102b; // 00400150: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h055: data = 32'h1440fff5; // 00400154: BNE, PC<=(REG[2] != REG[0])?PC+4+65525*4:PC+4;
      10'h056: data = 32'h00000000; // 00400158: SLL, REG[0]<=REG[0]<<0;
      10'h057: data = 32'h0810000d; // 0040015c: J, PC<=0x0010000d*4(=0x00400034);
      10'h058: data = 32'h00000000; // 00400160: SLL, REG[0]<=REG[0]<<0;
      10'h059: data = 32'hafc00014; // 00400164: SW, RAM[REG[30]+20]<=REG[0];
      10'h05a: data = 32'h08100062; // 00400168: J, PC<=0x00100062*4(=0x00400188);
      10'h05b: data = 32'h00000000; // 0040016c: SLL, REG[0]<=REG[0]<<0;
      10'h05c: data = 32'h0c100096; // 00400170: JAL, PC<=0x00100096*4(=0x00400258); REG[31]<=PC+4
      10'h05d: data = 32'h00000000; // 00400174: SLL, REG[0]<=REG[0]<<0;
      10'h05e: data = 32'h8fc20014; // 00400178: LW, REG[2]<=RAM[REG[30]+20];
      10'h05f: data = 32'h00000000; // 0040017c: SLL, REG[0]<=REG[0]<<0;
      10'h060: data = 32'h24420001; // 00400180: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h061: data = 32'hafc20014; // 00400184: SW, RAM[REG[30]+20]<=REG[2];
      10'h062: data = 32'h8fc20014; // 00400188: LW, REG[2]<=RAM[REG[30]+20];
      10'h063: data = 32'h8fc30010; // 0040018c: LW, REG[3]<=RAM[REG[30]+16];
      10'h064: data = 32'h00000000; // 00400190: SLL, REG[0]<=REG[0]<<0;
      10'h065: data = 32'h0043102b; // 00400194: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h066: data = 32'h1440fff5; // 00400198: BNE, PC<=(REG[2] != REG[0])?PC+4+65525*4:PC+4;
      10'h067: data = 32'h00000000; // 0040019c: SLL, REG[0]<=REG[0]<<0;
      10'h068: data = 32'h0810000d; // 004001a0: J, PC<=0x0010000d*4(=0x00400034);
      10'h069: data = 32'h00000000; // 004001a4: SLL, REG[0]<=REG[0]<<0;
      10'h06a: data = 32'h27bdffe8; // 004001a8: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h06b: data = 32'hafbf0014; // 004001ac: SW, RAM[REG[29]+20]<=REG[31];
      10'h06c: data = 32'hafbe0010; // 004001b0: SW, RAM[REG[29]+16]<=REG[30];
      10'h06d: data = 32'h03a0f021; // 004001b4: ADDU, REG[30]<=REG[29]+REG[0];
      10'h06e: data = 32'h24040008; // 004001b8: ADDIU, REG[4]<=REG[0]+8(=0x00000008);
      10'h06f: data = 32'h0c1000ac; // 004001bc: JAL, PC<=0x001000ac*4(=0x004002b0); REG[31]<=PC+4
      10'h070: data = 32'h00000000; // 004001c0: SLL, REG[0]<=REG[0]<<0;
      10'h071: data = 32'h24040004; // 004001c4: ADDIU, REG[4]<=REG[0]+4(=0x00000004);
      10'h072: data = 32'h0c1000ac; // 004001c8: JAL, PC<=0x001000ac*4(=0x004002b0); REG[31]<=PC+4
      10'h073: data = 32'h00000000; // 004001cc: SLL, REG[0]<=REG[0]<<0;
      10'h074: data = 32'h24040002; // 004001d0: ADDIU, REG[4]<=REG[0]+2(=0x00000002);
      10'h075: data = 32'h0c1000ac; // 004001d4: JAL, PC<=0x001000ac*4(=0x004002b0); REG[31]<=PC+4
      10'h076: data = 32'h00000000; // 004001d8: SLL, REG[0]<=REG[0]<<0;
      10'h077: data = 32'h24040001; // 004001dc: ADDIU, REG[4]<=REG[0]+1(=0x00000001);
      10'h078: data = 32'h0c1000ac; // 004001e0: JAL, PC<=0x001000ac*4(=0x004002b0); REG[31]<=PC+4
      10'h079: data = 32'h00000000; // 004001e4: SLL, REG[0]<=REG[0]<<0;
      10'h07a: data = 32'h03c0e821; // 004001e8: ADDU, REG[29]<=REG[30]+REG[0];
      10'h07b: data = 32'h8fbf0014; // 004001ec: LW, REG[31]<=RAM[REG[29]+20];
      10'h07c: data = 32'h8fbe0010; // 004001f0: LW, REG[30]<=RAM[REG[29]+16];
      10'h07d: data = 32'h27bd0018; // 004001f4: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h07e: data = 32'h03e00008; // 004001f8: JR, PC<=REG[31];
      10'h07f: data = 32'h00000000; // 004001fc: SLL, REG[0]<=REG[0]<<0;
      10'h080: data = 32'h27bdffe8; // 00400200: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h081: data = 32'hafbf0014; // 00400204: SW, RAM[REG[29]+20]<=REG[31];
      10'h082: data = 32'hafbe0010; // 00400208: SW, RAM[REG[29]+16]<=REG[30];
      10'h083: data = 32'h03a0f021; // 0040020c: ADDU, REG[30]<=REG[29]+REG[0];
      10'h084: data = 32'h24040008; // 00400210: ADDIU, REG[4]<=REG[0]+8(=0x00000008);
      10'h085: data = 32'h0c1000ac; // 00400214: JAL, PC<=0x001000ac*4(=0x004002b0); REG[31]<=PC+4
      10'h086: data = 32'h00000000; // 00400218: SLL, REG[0]<=REG[0]<<0;
      10'h087: data = 32'h24040001; // 0040021c: ADDIU, REG[4]<=REG[0]+1(=0x00000001);
      10'h088: data = 32'h0c1000ac; // 00400220: JAL, PC<=0x001000ac*4(=0x004002b0); REG[31]<=PC+4
      10'h089: data = 32'h00000000; // 00400224: SLL, REG[0]<=REG[0]<<0;
      10'h08a: data = 32'h24040002; // 00400228: ADDIU, REG[4]<=REG[0]+2(=0x00000002);
      10'h08b: data = 32'h0c1000ac; // 0040022c: JAL, PC<=0x001000ac*4(=0x004002b0); REG[31]<=PC+4
      10'h08c: data = 32'h00000000; // 00400230: SLL, REG[0]<=REG[0]<<0;
      10'h08d: data = 32'h24040004; // 00400234: ADDIU, REG[4]<=REG[0]+4(=0x00000004);
      10'h08e: data = 32'h0c1000ac; // 00400238: JAL, PC<=0x001000ac*4(=0x004002b0); REG[31]<=PC+4
      10'h08f: data = 32'h00000000; // 0040023c: SLL, REG[0]<=REG[0]<<0;
      10'h090: data = 32'h03c0e821; // 00400240: ADDU, REG[29]<=REG[30]+REG[0];
      10'h091: data = 32'h8fbf0014; // 00400244: LW, REG[31]<=RAM[REG[29]+20];
      10'h092: data = 32'h8fbe0010; // 00400248: LW, REG[30]<=RAM[REG[29]+16];
      10'h093: data = 32'h27bd0018; // 0040024c: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h094: data = 32'h03e00008; // 00400250: JR, PC<=REG[31];
      10'h095: data = 32'h00000000; // 00400254: SLL, REG[0]<=REG[0]<<0;
      10'h096: data = 32'h27bdffe8; // 00400258: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h097: data = 32'hafbf0014; // 0040025c: SW, RAM[REG[29]+20]<=REG[31];
      10'h098: data = 32'hafbe0010; // 00400260: SW, RAM[REG[29]+16]<=REG[30];
      10'h099: data = 32'h03a0f021; // 00400264: ADDU, REG[30]<=REG[29]+REG[0];
      10'h09a: data = 32'h24040008; // 00400268: ADDIU, REG[4]<=REG[0]+8(=0x00000008);
      10'h09b: data = 32'h0c1000ac; // 0040026c: JAL, PC<=0x001000ac*4(=0x004002b0); REG[31]<=PC+4
      10'h09c: data = 32'h00000000; // 00400270: SLL, REG[0]<=REG[0]<<0;
      10'h09d: data = 32'h24040008; // 00400274: ADDIU, REG[4]<=REG[0]+8(=0x00000008);
      10'h09e: data = 32'h0c1000ac; // 00400278: JAL, PC<=0x001000ac*4(=0x004002b0); REG[31]<=PC+4
      10'h09f: data = 32'h00000000; // 0040027c: SLL, REG[0]<=REG[0]<<0;
      10'h0a0: data = 32'h24040008; // 00400280: ADDIU, REG[4]<=REG[0]+8(=0x00000008);
      10'h0a1: data = 32'h0c1000ac; // 00400284: JAL, PC<=0x001000ac*4(=0x004002b0); REG[31]<=PC+4
      10'h0a2: data = 32'h00000000; // 00400288: SLL, REG[0]<=REG[0]<<0;
      10'h0a3: data = 32'h24040008; // 0040028c: ADDIU, REG[4]<=REG[0]+8(=0x00000008);
      10'h0a4: data = 32'h0c1000ac; // 00400290: JAL, PC<=0x001000ac*4(=0x004002b0); REG[31]<=PC+4
      10'h0a5: data = 32'h00000000; // 00400294: SLL, REG[0]<=REG[0]<<0;
      10'h0a6: data = 32'h03c0e821; // 00400298: ADDU, REG[29]<=REG[30]+REG[0];
      10'h0a7: data = 32'h8fbf0014; // 0040029c: LW, REG[31]<=RAM[REG[29]+20];
      10'h0a8: data = 32'h8fbe0010; // 004002a0: LW, REG[30]<=RAM[REG[29]+16];
      10'h0a9: data = 32'h27bd0018; // 004002a4: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h0aa: data = 32'h03e00008; // 004002a8: JR, PC<=REG[31];
      10'h0ab: data = 32'h00000000; // 004002ac: SLL, REG[0]<=REG[0]<<0;
      10'h0ac: data = 32'h27bdfff0; // 004002b0: ADDIU, REG[29]<=REG[29]+65520(=0x0000fff0);
      10'h0ad: data = 32'hafbe0008; // 004002b4: SW, RAM[REG[29]+8]<=REG[30];
      10'h0ae: data = 32'h03a0f021; // 004002b8: ADDU, REG[30]<=REG[29]+REG[0];
      10'h0af: data = 32'hafc40010; // 004002bc: SW, RAM[REG[30]+16]<=REG[4];
      10'h0b0: data = 32'h24030320; // 004002c0: ADDIU, REG[3]<=REG[0]+800(=0x00000320);
      10'h0b1: data = 32'h8fc20010; // 004002c4: LW, REG[2]<=RAM[REG[30]+16];
      10'h0b2: data = 32'h00000000; // 004002c8: SLL, REG[0]<=REG[0]<<0;
      10'h0b3: data = 32'hac620000; // 004002cc: SW, RAM[REG[3]+0]<=REG[2];
      10'h0b4: data = 32'h03c0e821; // 004002d0: ADDU, REG[29]<=REG[30]+REG[0];
      10'h0b5: data = 32'h8fbe0008; // 004002d4: LW, REG[30]<=RAM[REG[29]+8];
      10'h0b6: data = 32'h27bd0010; // 004002d8: ADDIU, REG[29]<=REG[29]+16(=0x00000010);
      10'h0b7: data = 32'h03e00008; // 004002dc: JR, PC<=REG[31];
      10'h0b8: data = 32'h00000000; // 004002e0: SLL, REG[0]<=REG[0]<<0;
      10'h0b9: data = 32'h27bdfff8; // 004002e4: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h0ba: data = 32'hafbe0000; // 004002e8: SW, RAM[REG[29]+0]<=REG[30];
      10'h0bb: data = 32'h03a0f021; // 004002ec: ADDU, REG[30]<=REG[29]+REG[0];
      10'h0bc: data = 32'hafc40008; // 004002f0: SW, RAM[REG[30]+8]<=REG[4];
      10'h0bd: data = 32'h24020308; // 004002f4: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h0be: data = 32'hac400000; // 004002f8: SW, RAM[REG[2]+0]<=REG[0];
      10'h0bf: data = 32'h2403030c; // 004002fc: ADDIU, REG[3]<=REG[0]+780(=0x0000030c);
      10'h0c0: data = 32'h24020001; // 00400300: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0c1: data = 32'hac620000; // 00400304: SW, RAM[REG[3]+0]<=REG[2];
      10'h0c2: data = 32'h24030308; // 00400308: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h0c3: data = 32'h24020001; // 0040030c: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0c4: data = 32'hac620000; // 00400310: SW, RAM[REG[3]+0]<=REG[2];
      10'h0c5: data = 32'h24020308; // 00400314: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h0c6: data = 32'hac400000; // 00400318: SW, RAM[REG[2]+0]<=REG[0];
      10'h0c7: data = 32'h24030308; // 0040031c: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h0c8: data = 32'h24020001; // 00400320: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0c9: data = 32'hac620000; // 00400324: SW, RAM[REG[3]+0]<=REG[2];
      10'h0ca: data = 32'h081000d1; // 00400328: J, PC<=0x001000d1*4(=0x00400344);
      10'h0cb: data = 32'h00000000; // 0040032c: SLL, REG[0]<=REG[0]<<0;
      10'h0cc: data = 32'h24020308; // 00400330: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h0cd: data = 32'hac400000; // 00400334: SW, RAM[REG[2]+0]<=REG[0];
      10'h0ce: data = 32'h24030308; // 00400338: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h0cf: data = 32'h24020001; // 0040033c: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0d0: data = 32'hac620000; // 00400340: SW, RAM[REG[3]+0]<=REG[2];
      10'h0d1: data = 32'h24020310; // 00400344: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h0d2: data = 32'h8c430000; // 00400348: LW, REG[3]<=RAM[REG[2]+0];
      10'h0d3: data = 32'h2402ffff; // 0040034c: ADDIU, REG[2]<=REG[0]+65535(=0x0000ffff);
      10'h0d4: data = 32'h1062fff7; // 00400350: BEQ, PC<=(REG[3] == REG[2])?PC+4+65527*4:PC+4;
      10'h0d5: data = 32'h00000000; // 00400354: SLL, REG[0]<=REG[0]<<0;
      10'h0d6: data = 32'h0810017f; // 00400358: J, PC<=0x0010017f*4(=0x004005fc);
      10'h0d7: data = 32'h00000000; // 0040035c: SLL, REG[0]<=REG[0]<<0;
      10'h0d8: data = 32'h8fc20008; // 00400360: LW, REG[2]<=RAM[REG[30]+8];
      10'h0d9: data = 32'h00000000; // 00400364: SLL, REG[0]<=REG[0]<<0;
      10'h0da: data = 32'h8c420000; // 00400368: LW, REG[2]<=RAM[REG[2]+0];
      10'h0db: data = 32'h00000000; // 0040036c: SLL, REG[0]<=REG[0]<<0;
      10'h0dc: data = 32'h10400012; // 00400370: BEQ, PC<=(REG[2] == REG[0])?PC+4+18*4:PC+4;
      10'h0dd: data = 32'h00000000; // 00400374: SLL, REG[0]<=REG[0]<<0;
      10'h0de: data = 32'h8fc20008; // 00400378: LW, REG[2]<=RAM[REG[30]+8];
      10'h0df: data = 32'h00000000; // 0040037c: SLL, REG[0]<=REG[0]<<0;
      10'h0e0: data = 32'h8c420000; // 00400380: LW, REG[2]<=RAM[REG[2]+0];
      10'h0e1: data = 32'h00000000; // 00400384: SLL, REG[0]<=REG[0]<<0;
      10'h0e2: data = 32'h2c42001b; // 00400388: SLTIU, REG[2]<=(REG[2]<27(=0x0000001b))?1:0;
      10'h0e3: data = 32'h1040000b; // 0040038c: BEQ, PC<=(REG[2] == REG[0])?PC+4+11*4:PC+4;
      10'h0e4: data = 32'h00000000; // 00400390: SLL, REG[0]<=REG[0]<<0;
      10'h0e5: data = 32'h8fc20008; // 00400394: LW, REG[2]<=RAM[REG[30]+8];
      10'h0e6: data = 32'h00000000; // 00400398: SLL, REG[0]<=REG[0]<<0;
      10'h0e7: data = 32'h8c420000; // 0040039c: LW, REG[2]<=RAM[REG[2]+0];
      10'h0e8: data = 32'h00000000; // 004003a0: SLL, REG[0]<=REG[0]<<0;
      10'h0e9: data = 32'h24430040; // 004003a4: ADDIU, REG[3]<=REG[2]+64(=0x00000040);
      10'h0ea: data = 32'h8fc20008; // 004003a8: LW, REG[2]<=RAM[REG[30]+8];
      10'h0eb: data = 32'h00000000; // 004003ac: SLL, REG[0]<=REG[0]<<0;
      10'h0ec: data = 32'hac430000; // 004003b0: SW, RAM[REG[2]+0]<=REG[3];
      10'h0ed: data = 32'h08100176; // 004003b4: J, PC<=0x00100176*4(=0x004005d8);
      10'h0ee: data = 32'h00000000; // 004003b8: SLL, REG[0]<=REG[0]<<0;
      10'h0ef: data = 32'h8fc20008; // 004003bc: LW, REG[2]<=RAM[REG[30]+8];
      10'h0f0: data = 32'h00000000; // 004003c0: SLL, REG[0]<=REG[0]<<0;
      10'h0f1: data = 32'h8c420000; // 004003c4: LW, REG[2]<=RAM[REG[2]+0];
      10'h0f2: data = 32'h00000000; // 004003c8: SLL, REG[0]<=REG[0]<<0;
      10'h0f3: data = 32'h2c420030; // 004003cc: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h0f4: data = 32'h14400010; // 004003d0: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h0f5: data = 32'h00000000; // 004003d4: SLL, REG[0]<=REG[0]<<0;
      10'h0f6: data = 32'h8fc20008; // 004003d8: LW, REG[2]<=RAM[REG[30]+8];
      10'h0f7: data = 32'h00000000; // 004003dc: SLL, REG[0]<=REG[0]<<0;
      10'h0f8: data = 32'h8c420000; // 004003e0: LW, REG[2]<=RAM[REG[2]+0];
      10'h0f9: data = 32'h00000000; // 004003e4: SLL, REG[0]<=REG[0]<<0;
      10'h0fa: data = 32'h2c42003a; // 004003e8: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h0fb: data = 32'h10400009; // 004003ec: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h0fc: data = 32'h00000000; // 004003f0: SLL, REG[0]<=REG[0]<<0;
      10'h0fd: data = 32'h8fc20008; // 004003f4: LW, REG[2]<=RAM[REG[30]+8];
      10'h0fe: data = 32'h00000000; // 004003f8: SLL, REG[0]<=REG[0]<<0;
      10'h0ff: data = 32'h8c430000; // 004003fc: LW, REG[3]<=RAM[REG[2]+0];
      10'h100: data = 32'h8fc20008; // 00400400: LW, REG[2]<=RAM[REG[30]+8];
      10'h101: data = 32'h00000000; // 00400404: SLL, REG[0]<=REG[0]<<0;
      10'h102: data = 32'hac430000; // 00400408: SW, RAM[REG[2]+0]<=REG[3];
      10'h103: data = 32'h08100176; // 0040040c: J, PC<=0x00100176*4(=0x004005d8);
      10'h104: data = 32'h00000000; // 00400410: SLL, REG[0]<=REG[0]<<0;
      10'h105: data = 32'h8fc20008; // 00400414: LW, REG[2]<=RAM[REG[30]+8];
      10'h106: data = 32'h00000000; // 00400418: SLL, REG[0]<=REG[0]<<0;
      10'h107: data = 32'h8c420000; // 0040041c: LW, REG[2]<=RAM[REG[2]+0];
      10'h108: data = 32'h00000000; // 00400420: SLL, REG[0]<=REG[0]<<0;
      10'h109: data = 32'h14400006; // 00400424: BNE, PC<=(REG[2] != REG[0])?PC+4+6*4:PC+4;
      10'h10a: data = 32'h00000000; // 00400428: SLL, REG[0]<=REG[0]<<0;
      10'h10b: data = 32'h8fc30008; // 0040042c: LW, REG[3]<=RAM[REG[30]+8];
      10'h10c: data = 32'h24020040; // 00400430: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h10d: data = 32'hac620000; // 00400434: SW, RAM[REG[3]+0]<=REG[2];
      10'h10e: data = 32'h08100176; // 00400438: J, PC<=0x00100176*4(=0x004005d8);
      10'h10f: data = 32'h00000000; // 0040043c: SLL, REG[0]<=REG[0]<<0;
      10'h110: data = 32'h8fc20008; // 00400440: LW, REG[2]<=RAM[REG[30]+8];
      10'h111: data = 32'h00000000; // 00400444: SLL, REG[0]<=REG[0]<<0;
      10'h112: data = 32'h8c430000; // 00400448: LW, REG[3]<=RAM[REG[2]+0];
      10'h113: data = 32'h2402001b; // 0040044c: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h114: data = 32'h14620006; // 00400450: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h115: data = 32'h00000000; // 00400454: SLL, REG[0]<=REG[0]<<0;
      10'h116: data = 32'h8fc30008; // 00400458: LW, REG[3]<=RAM[REG[30]+8];
      10'h117: data = 32'h2402005b; // 0040045c: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h118: data = 32'hac620000; // 00400460: SW, RAM[REG[3]+0]<=REG[2];
      10'h119: data = 32'h08100176; // 00400464: J, PC<=0x00100176*4(=0x004005d8);
      10'h11a: data = 32'h00000000; // 00400468: SLL, REG[0]<=REG[0]<<0;
      10'h11b: data = 32'h8fc20008; // 0040046c: LW, REG[2]<=RAM[REG[30]+8];
      10'h11c: data = 32'h00000000; // 00400470: SLL, REG[0]<=REG[0]<<0;
      10'h11d: data = 32'h8c430000; // 00400474: LW, REG[3]<=RAM[REG[2]+0];
      10'h11e: data = 32'h2402001d; // 00400478: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h11f: data = 32'h14620006; // 0040047c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h120: data = 32'h00000000; // 00400480: SLL, REG[0]<=REG[0]<<0;
      10'h121: data = 32'h8fc30008; // 00400484: LW, REG[3]<=RAM[REG[30]+8];
      10'h122: data = 32'h2402005d; // 00400488: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h123: data = 32'hac620000; // 0040048c: SW, RAM[REG[3]+0]<=REG[2];
      10'h124: data = 32'h08100176; // 00400490: J, PC<=0x00100176*4(=0x004005d8);
      10'h125: data = 32'h00000000; // 00400494: SLL, REG[0]<=REG[0]<<0;
      10'h126: data = 32'h8fc20008; // 00400498: LW, REG[2]<=RAM[REG[30]+8];
      10'h127: data = 32'h00000000; // 0040049c: SLL, REG[0]<=REG[0]<<0;
      10'h128: data = 32'h8c420000; // 004004a0: LW, REG[2]<=RAM[REG[2]+0];
      10'h129: data = 32'h00000000; // 004004a4: SLL, REG[0]<=REG[0]<<0;
      10'h12a: data = 32'h2c420020; // 004004a8: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h12b: data = 32'h14400010; // 004004ac: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h12c: data = 32'h00000000; // 004004b0: SLL, REG[0]<=REG[0]<<0;
      10'h12d: data = 32'h8fc20008; // 004004b4: LW, REG[2]<=RAM[REG[30]+8];
      10'h12e: data = 32'h00000000; // 004004b8: SLL, REG[0]<=REG[0]<<0;
      10'h12f: data = 32'h8c420000; // 004004bc: LW, REG[2]<=RAM[REG[2]+0];
      10'h130: data = 32'h00000000; // 004004c0: SLL, REG[0]<=REG[0]<<0;
      10'h131: data = 32'h2c420030; // 004004c4: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h132: data = 32'h10400009; // 004004c8: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h133: data = 32'h00000000; // 004004cc: SLL, REG[0]<=REG[0]<<0;
      10'h134: data = 32'h8fc20008; // 004004d0: LW, REG[2]<=RAM[REG[30]+8];
      10'h135: data = 32'h00000000; // 004004d4: SLL, REG[0]<=REG[0]<<0;
      10'h136: data = 32'h8c430000; // 004004d8: LW, REG[3]<=RAM[REG[2]+0];
      10'h137: data = 32'h8fc20008; // 004004dc: LW, REG[2]<=RAM[REG[30]+8];
      10'h138: data = 32'h00000000; // 004004e0: SLL, REG[0]<=REG[0]<<0;
      10'h139: data = 32'hac430000; // 004004e4: SW, RAM[REG[2]+0]<=REG[3];
      10'h13a: data = 32'h08100176; // 004004e8: J, PC<=0x00100176*4(=0x004005d8);
      10'h13b: data = 32'h00000000; // 004004ec: SLL, REG[0]<=REG[0]<<0;
      10'h13c: data = 32'h8fc20008; // 004004f0: LW, REG[2]<=RAM[REG[30]+8];
      10'h13d: data = 32'h00000000; // 004004f4: SLL, REG[0]<=REG[0]<<0;
      10'h13e: data = 32'h8c430000; // 004004f8: LW, REG[3]<=RAM[REG[2]+0];
      10'h13f: data = 32'h2402003a; // 004004fc: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h140: data = 32'h14620006; // 00400500: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h141: data = 32'h00000000; // 00400504: SLL, REG[0]<=REG[0]<<0;
      10'h142: data = 32'h8fc30008; // 00400508: LW, REG[3]<=RAM[REG[30]+8];
      10'h143: data = 32'h2402003f; // 0040050c: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h144: data = 32'hac620000; // 00400510: SW, RAM[REG[3]+0]<=REG[2];
      10'h145: data = 32'h08100176; // 00400514: J, PC<=0x00100176*4(=0x004005d8);
      10'h146: data = 32'h00000000; // 00400518: SLL, REG[0]<=REG[0]<<0;
      10'h147: data = 32'h8fc20008; // 0040051c: LW, REG[2]<=RAM[REG[30]+8];
      10'h148: data = 32'h00000000; // 00400520: SLL, REG[0]<=REG[0]<<0;
      10'h149: data = 32'h8c430000; // 00400524: LW, REG[3]<=RAM[REG[2]+0];
      10'h14a: data = 32'h2402003b; // 00400528: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h14b: data = 32'h14620006; // 0040052c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h14c: data = 32'h00000000; // 00400530: SLL, REG[0]<=REG[0]<<0;
      10'h14d: data = 32'h8fc30008; // 00400534: LW, REG[3]<=RAM[REG[30]+8];
      10'h14e: data = 32'h2402003d; // 00400538: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h14f: data = 32'hac620000; // 0040053c: SW, RAM[REG[3]+0]<=REG[2];
      10'h150: data = 32'h08100176; // 00400540: J, PC<=0x00100176*4(=0x004005d8);
      10'h151: data = 32'h00000000; // 00400544: SLL, REG[0]<=REG[0]<<0;
      10'h152: data = 32'h8fc20008; // 00400548: LW, REG[2]<=RAM[REG[30]+8];
      10'h153: data = 32'h00000000; // 0040054c: SLL, REG[0]<=REG[0]<<0;
      10'h154: data = 32'h8c430000; // 00400550: LW, REG[3]<=RAM[REG[2]+0];
      10'h155: data = 32'h2402003c; // 00400554: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h156: data = 32'h14620006; // 00400558: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h157: data = 32'h00000000; // 0040055c: SLL, REG[0]<=REG[0]<<0;
      10'h158: data = 32'h8fc30008; // 00400560: LW, REG[3]<=RAM[REG[30]+8];
      10'h159: data = 32'h2402003b; // 00400564: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h15a: data = 32'hac620000; // 00400568: SW, RAM[REG[3]+0]<=REG[2];
      10'h15b: data = 32'h08100176; // 0040056c: J, PC<=0x00100176*4(=0x004005d8);
      10'h15c: data = 32'h00000000; // 00400570: SLL, REG[0]<=REG[0]<<0;
      10'h15d: data = 32'h8fc20008; // 00400574: LW, REG[2]<=RAM[REG[30]+8];
      10'h15e: data = 32'h00000000; // 00400578: SLL, REG[0]<=REG[0]<<0;
      10'h15f: data = 32'h8c430000; // 0040057c: LW, REG[3]<=RAM[REG[2]+0];
      10'h160: data = 32'h2402003d; // 00400580: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h161: data = 32'h14620006; // 00400584: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h162: data = 32'h00000000; // 00400588: SLL, REG[0]<=REG[0]<<0;
      10'h163: data = 32'h8fc30008; // 0040058c: LW, REG[3]<=RAM[REG[30]+8];
      10'h164: data = 32'h2402003a; // 00400590: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h165: data = 32'hac620000; // 00400594: SW, RAM[REG[3]+0]<=REG[2];
      10'h166: data = 32'h08100176; // 00400598: J, PC<=0x00100176*4(=0x004005d8);
      10'h167: data = 32'h00000000; // 0040059c: SLL, REG[0]<=REG[0]<<0;
      10'h168: data = 32'h8fc20008; // 004005a0: LW, REG[2]<=RAM[REG[30]+8];
      10'h169: data = 32'h00000000; // 004005a4: SLL, REG[0]<=REG[0]<<0;
      10'h16a: data = 32'h8c430000; // 004005a8: LW, REG[3]<=RAM[REG[2]+0];
      10'h16b: data = 32'h2402003e; // 004005ac: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h16c: data = 32'h14620006; // 004005b0: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h16d: data = 32'h00000000; // 004005b4: SLL, REG[0]<=REG[0]<<0;
      10'h16e: data = 32'h8fc30008; // 004005b8: LW, REG[3]<=RAM[REG[30]+8];
      10'h16f: data = 32'h2402000a; // 004005bc: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h170: data = 32'hac620000; // 004005c0: SW, RAM[REG[3]+0]<=REG[2];
      10'h171: data = 32'h08100176; // 004005c4: J, PC<=0x00100176*4(=0x004005d8);
      10'h172: data = 32'h00000000; // 004005c8: SLL, REG[0]<=REG[0]<<0;
      10'h173: data = 32'h8fc30008; // 004005cc: LW, REG[3]<=RAM[REG[30]+8];
      10'h174: data = 32'h24020040; // 004005d0: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h175: data = 32'hac620000; // 004005d4: SW, RAM[REG[3]+0]<=REG[2];
      10'h176: data = 32'h24020308; // 004005d8: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h177: data = 32'hac400000; // 004005dc: SW, RAM[REG[2]+0]<=REG[0];
      10'h178: data = 32'h24030308; // 004005e0: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h179: data = 32'h24020001; // 004005e4: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h17a: data = 32'hac620000; // 004005e8: SW, RAM[REG[3]+0]<=REG[2];
      10'h17b: data = 32'h8fc20008; // 004005ec: LW, REG[2]<=RAM[REG[30]+8];
      10'h17c: data = 32'h00000000; // 004005f0: SLL, REG[0]<=REG[0]<<0;
      10'h17d: data = 32'h24420004; // 004005f4: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h17e: data = 32'hafc20008; // 004005f8: SW, RAM[REG[30]+8]<=REG[2];
      10'h17f: data = 32'h24020310; // 004005fc: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h180: data = 32'h8c430000; // 00400600: LW, REG[3]<=RAM[REG[2]+0];
      10'h181: data = 32'h8fc20008; // 00400604: LW, REG[2]<=RAM[REG[30]+8];
      10'h182: data = 32'h00000000; // 00400608: SLL, REG[0]<=REG[0]<<0;
      10'h183: data = 32'hac430000; // 0040060c: SW, RAM[REG[2]+0]<=REG[3];
      10'h184: data = 32'h8fc20008; // 00400610: LW, REG[2]<=RAM[REG[30]+8];
      10'h185: data = 32'h00000000; // 00400614: SLL, REG[0]<=REG[0]<<0;
      10'h186: data = 32'h8c430000; // 00400618: LW, REG[3]<=RAM[REG[2]+0];
      10'h187: data = 32'h2402003e; // 0040061c: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h188: data = 32'h1462ff4f; // 00400620: BNE, PC<=(REG[3] != REG[2])?PC+4+65359*4:PC+4;
      10'h189: data = 32'h00000000; // 00400624: SLL, REG[0]<=REG[0]<<0;
      10'h18a: data = 32'h8fc20008; // 00400628: LW, REG[2]<=RAM[REG[30]+8];
      10'h18b: data = 32'h00000000; // 0040062c: SLL, REG[0]<=REG[0]<<0;
      10'h18c: data = 32'hac400000; // 00400630: SW, RAM[REG[2]+0]<=REG[0];
      10'h18d: data = 32'h24020308; // 00400634: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h18e: data = 32'hac400000; // 00400638: SW, RAM[REG[2]+0]<=REG[0];
      10'h18f: data = 32'h2402030c; // 0040063c: ADDIU, REG[2]<=REG[0]+780(=0x0000030c);
      10'h190: data = 32'hac400000; // 00400640: SW, RAM[REG[2]+0]<=REG[0];
      10'h191: data = 32'h24030308; // 00400644: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h192: data = 32'h24020001; // 00400648: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h193: data = 32'hac620000; // 0040064c: SW, RAM[REG[3]+0]<=REG[2];
      10'h194: data = 32'h24020308; // 00400650: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h195: data = 32'hac400000; // 00400654: SW, RAM[REG[2]+0]<=REG[0];
      10'h196: data = 32'h03c0e821; // 00400658: ADDU, REG[29]<=REG[30]+REG[0];
      10'h197: data = 32'h8fbe0000; // 0040065c: LW, REG[30]<=RAM[REG[29]+0];
      10'h198: data = 32'h27bd0008; // 00400660: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h199: data = 32'h03e00008; // 00400664: JR, PC<=REG[31];
      10'h19a: data = 32'h00000000; // 00400668: SLL, REG[0]<=REG[0]<<0;
      10'h19b: data = 32'h27bdffe8; // 0040066c: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h19c: data = 32'hafbe0010; // 00400670: SW, RAM[REG[29]+16]<=REG[30];
      10'h19d: data = 32'h03a0f021; // 00400674: ADDU, REG[30]<=REG[29]+REG[0];
      10'h19e: data = 32'hafc40018; // 00400678: SW, RAM[REG[30]+24]<=REG[4];
      10'h19f: data = 32'h8fc20018; // 0040067c: LW, REG[2]<=RAM[REG[30]+24];
      10'h1a0: data = 32'h00000000; // 00400680: SLL, REG[0]<=REG[0]<<0;
      10'h1a1: data = 32'hafc20008; // 00400684: SW, RAM[REG[30]+8]<=REG[2];
      10'h1a2: data = 32'hafc00004; // 00400688: SW, RAM[REG[30]+4]<=REG[0];
      10'h1a3: data = 32'h081001ad; // 0040068c: J, PC<=0x001001ad*4(=0x004006b4);
      10'h1a4: data = 32'h00000000; // 00400690: SLL, REG[0]<=REG[0]<<0;
      10'h1a5: data = 32'h8fc20008; // 00400694: LW, REG[2]<=RAM[REG[30]+8];
      10'h1a6: data = 32'h00000000; // 00400698: SLL, REG[0]<=REG[0]<<0;
      10'h1a7: data = 32'h24420004; // 0040069c: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h1a8: data = 32'hafc20008; // 004006a0: SW, RAM[REG[30]+8]<=REG[2];
      10'h1a9: data = 32'h8fc20004; // 004006a4: LW, REG[2]<=RAM[REG[30]+4];
      10'h1aa: data = 32'h00000000; // 004006a8: SLL, REG[0]<=REG[0]<<0;
      10'h1ab: data = 32'h24420001; // 004006ac: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h1ac: data = 32'hafc20004; // 004006b0: SW, RAM[REG[30]+4]<=REG[2];
      10'h1ad: data = 32'h8fc20008; // 004006b4: LW, REG[2]<=RAM[REG[30]+8];
      10'h1ae: data = 32'h00000000; // 004006b8: SLL, REG[0]<=REG[0]<<0;
      10'h1af: data = 32'h8c420000; // 004006bc: LW, REG[2]<=RAM[REG[2]+0];
      10'h1b0: data = 32'h00000000; // 004006c0: SLL, REG[0]<=REG[0]<<0;
      10'h1b1: data = 32'h1440fff3; // 004006c4: BNE, PC<=(REG[2] != REG[0])?PC+4+65523*4:PC+4;
      10'h1b2: data = 32'h00000000; // 004006c8: SLL, REG[0]<=REG[0]<<0;
      10'h1b3: data = 32'hafc00000; // 004006cc: SW, RAM[REG[30]+0]<=REG[0];
      10'h1b4: data = 32'h8fc20018; // 004006d0: LW, REG[2]<=RAM[REG[30]+24];
      10'h1b5: data = 32'h00000000; // 004006d4: SLL, REG[0]<=REG[0]<<0;
      10'h1b6: data = 32'hafc20008; // 004006d8: SW, RAM[REG[30]+8]<=REG[2];
      10'h1b7: data = 32'h8fc30004; // 004006dc: LW, REG[3]<=RAM[REG[30]+4];
      10'h1b8: data = 32'h24020001; // 004006e0: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h1b9: data = 32'h14620009; // 004006e4: BNE, PC<=(REG[3] != REG[2])?PC+4+9*4:PC+4;
      10'h1ba: data = 32'h00000000; // 004006e8: SLL, REG[0]<=REG[0]<<0;
      10'h1bb: data = 32'h8fc20008; // 004006ec: LW, REG[2]<=RAM[REG[30]+8];
      10'h1bc: data = 32'h00000000; // 004006f0: SLL, REG[0]<=REG[0]<<0;
      10'h1bd: data = 32'h8c420000; // 004006f4: LW, REG[2]<=RAM[REG[2]+0];
      10'h1be: data = 32'h00000000; // 004006f8: SLL, REG[0]<=REG[0]<<0;
      10'h1bf: data = 32'h2442ffd0; // 004006fc: ADDIU, REG[2]<=REG[2]+65488(=0x0000ffd0);
      10'h1c0: data = 32'hafc20000; // 00400700: SW, RAM[REG[30]+0]<=REG[2];
      10'h1c1: data = 32'h08100228; // 00400704: J, PC<=0x00100228*4(=0x004008a0);
      10'h1c2: data = 32'h00000000; // 00400708: SLL, REG[0]<=REG[0]<<0;
      10'h1c3: data = 32'h8fc30004; // 0040070c: LW, REG[3]<=RAM[REG[30]+4];
      10'h1c4: data = 32'h24020002; // 00400710: ADDIU, REG[2]<=REG[0]+2(=0x00000002);
      10'h1c5: data = 32'h14620024; // 00400714: BNE, PC<=(REG[3] != REG[2])?PC+4+36*4:PC+4;
      10'h1c6: data = 32'h00000000; // 00400718: SLL, REG[0]<=REG[0]<<0;
      10'h1c7: data = 32'hafc00004; // 0040071c: SW, RAM[REG[30]+4]<=REG[0];
      10'h1c8: data = 32'h081001d2; // 00400720: J, PC<=0x001001d2*4(=0x00400748);
      10'h1c9: data = 32'h00000000; // 00400724: SLL, REG[0]<=REG[0]<<0;
      10'h1ca: data = 32'h8fc20000; // 00400728: LW, REG[2]<=RAM[REG[30]+0];
      10'h1cb: data = 32'h00000000; // 0040072c: SLL, REG[0]<=REG[0]<<0;
      10'h1cc: data = 32'h2442000a; // 00400730: ADDIU, REG[2]<=REG[2]+10(=0x0000000a);
      10'h1cd: data = 32'hafc20000; // 00400734: SW, RAM[REG[30]+0]<=REG[2];
      10'h1ce: data = 32'h8fc20004; // 00400738: LW, REG[2]<=RAM[REG[30]+4];
      10'h1cf: data = 32'h00000000; // 0040073c: SLL, REG[0]<=REG[0]<<0;
      10'h1d0: data = 32'h24420001; // 00400740: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h1d1: data = 32'hafc20004; // 00400744: SW, RAM[REG[30]+4]<=REG[2];
      10'h1d2: data = 32'h8fc20008; // 00400748: LW, REG[2]<=RAM[REG[30]+8];
      10'h1d3: data = 32'h00000000; // 0040074c: SLL, REG[0]<=REG[0]<<0;
      10'h1d4: data = 32'h8c420000; // 00400750: LW, REG[2]<=RAM[REG[2]+0];
      10'h1d5: data = 32'h00000000; // 00400754: SLL, REG[0]<=REG[0]<<0;
      10'h1d6: data = 32'h2443ffd0; // 00400758: ADDIU, REG[3]<=REG[2]+65488(=0x0000ffd0);
      10'h1d7: data = 32'h8fc20004; // 0040075c: LW, REG[2]<=RAM[REG[30]+4];
      10'h1d8: data = 32'h00000000; // 00400760: SLL, REG[0]<=REG[0]<<0;
      10'h1d9: data = 32'h0043102b; // 00400764: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h1da: data = 32'h1440ffef; // 00400768: BNE, PC<=(REG[2] != REG[0])?PC+4+65519*4:PC+4;
      10'h1db: data = 32'h00000000; // 0040076c: SLL, REG[0]<=REG[0]<<0;
      10'h1dc: data = 32'h8fc20008; // 00400770: LW, REG[2]<=RAM[REG[30]+8];
      10'h1dd: data = 32'h00000000; // 00400774: SLL, REG[0]<=REG[0]<<0;
      10'h1de: data = 32'h24420004; // 00400778: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h1df: data = 32'hafc20008; // 0040077c: SW, RAM[REG[30]+8]<=REG[2];
      10'h1e0: data = 32'h8fc20008; // 00400780: LW, REG[2]<=RAM[REG[30]+8];
      10'h1e1: data = 32'h00000000; // 00400784: SLL, REG[0]<=REG[0]<<0;
      10'h1e2: data = 32'h8c430000; // 00400788: LW, REG[3]<=RAM[REG[2]+0];
      10'h1e3: data = 32'h8fc20000; // 0040078c: LW, REG[2]<=RAM[REG[30]+0];
      10'h1e4: data = 32'h00000000; // 00400790: SLL, REG[0]<=REG[0]<<0;
      10'h1e5: data = 32'h00621021; // 00400794: ADDU, REG[2]<=REG[3]+REG[2];
      10'h1e6: data = 32'h2442ffd0; // 00400798: ADDIU, REG[2]<=REG[2]+65488(=0x0000ffd0);
      10'h1e7: data = 32'hafc20000; // 0040079c: SW, RAM[REG[30]+0]<=REG[2];
      10'h1e8: data = 32'h08100228; // 004007a0: J, PC<=0x00100228*4(=0x004008a0);
      10'h1e9: data = 32'h00000000; // 004007a4: SLL, REG[0]<=REG[0]<<0;
      10'h1ea: data = 32'h8fc30004; // 004007a8: LW, REG[3]<=RAM[REG[30]+4];
      10'h1eb: data = 32'h24020003; // 004007ac: ADDIU, REG[2]<=REG[0]+3(=0x00000003);
      10'h1ec: data = 32'h1462003b; // 004007b0: BNE, PC<=(REG[3] != REG[2])?PC+4+59*4:PC+4;
      10'h1ed: data = 32'h00000000; // 004007b4: SLL, REG[0]<=REG[0]<<0;
      10'h1ee: data = 32'hafc00004; // 004007b8: SW, RAM[REG[30]+4]<=REG[0];
      10'h1ef: data = 32'h081001f9; // 004007bc: J, PC<=0x001001f9*4(=0x004007e4);
      10'h1f0: data = 32'h00000000; // 004007c0: SLL, REG[0]<=REG[0]<<0;
      10'h1f1: data = 32'h8fc20000; // 004007c4: LW, REG[2]<=RAM[REG[30]+0];
      10'h1f2: data = 32'h00000000; // 004007c8: SLL, REG[0]<=REG[0]<<0;
      10'h1f3: data = 32'h24420064; // 004007cc: ADDIU, REG[2]<=REG[2]+100(=0x00000064);
      10'h1f4: data = 32'hafc20000; // 004007d0: SW, RAM[REG[30]+0]<=REG[2];
      10'h1f5: data = 32'h8fc20004; // 004007d4: LW, REG[2]<=RAM[REG[30]+4];
      10'h1f6: data = 32'h00000000; // 004007d8: SLL, REG[0]<=REG[0]<<0;
      10'h1f7: data = 32'h24420001; // 004007dc: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h1f8: data = 32'hafc20004; // 004007e0: SW, RAM[REG[30]+4]<=REG[2];
      10'h1f9: data = 32'h8fc20008; // 004007e4: LW, REG[2]<=RAM[REG[30]+8];
      10'h1fa: data = 32'h00000000; // 004007e8: SLL, REG[0]<=REG[0]<<0;
      10'h1fb: data = 32'h8c420000; // 004007ec: LW, REG[2]<=RAM[REG[2]+0];
      10'h1fc: data = 32'h00000000; // 004007f0: SLL, REG[0]<=REG[0]<<0;
      10'h1fd: data = 32'h2443ffd0; // 004007f4: ADDIU, REG[3]<=REG[2]+65488(=0x0000ffd0);
      10'h1fe: data = 32'h8fc20004; // 004007f8: LW, REG[2]<=RAM[REG[30]+4];
      10'h1ff: data = 32'h00000000; // 004007fc: SLL, REG[0]<=REG[0]<<0;
      10'h200: data = 32'h0043102b; // 00400800: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h201: data = 32'h1440ffef; // 00400804: BNE, PC<=(REG[2] != REG[0])?PC+4+65519*4:PC+4;
      10'h202: data = 32'h00000000; // 00400808: SLL, REG[0]<=REG[0]<<0;
      10'h203: data = 32'h8fc20008; // 0040080c: LW, REG[2]<=RAM[REG[30]+8];
      10'h204: data = 32'h00000000; // 00400810: SLL, REG[0]<=REG[0]<<0;
      10'h205: data = 32'h24420004; // 00400814: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h206: data = 32'hafc20008; // 00400818: SW, RAM[REG[30]+8]<=REG[2];
      10'h207: data = 32'hafc00004; // 0040081c: SW, RAM[REG[30]+4]<=REG[0];
      10'h208: data = 32'h08100212; // 00400820: J, PC<=0x00100212*4(=0x00400848);
      10'h209: data = 32'h00000000; // 00400824: SLL, REG[0]<=REG[0]<<0;
      10'h20a: data = 32'h8fc20000; // 00400828: LW, REG[2]<=RAM[REG[30]+0];
      10'h20b: data = 32'h00000000; // 0040082c: SLL, REG[0]<=REG[0]<<0;
      10'h20c: data = 32'h2442000a; // 00400830: ADDIU, REG[2]<=REG[2]+10(=0x0000000a);
      10'h20d: data = 32'hafc20000; // 00400834: SW, RAM[REG[30]+0]<=REG[2];
      10'h20e: data = 32'h8fc20004; // 00400838: LW, REG[2]<=RAM[REG[30]+4];
      10'h20f: data = 32'h00000000; // 0040083c: SLL, REG[0]<=REG[0]<<0;
      10'h210: data = 32'h24420001; // 00400840: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h211: data = 32'hafc20004; // 00400844: SW, RAM[REG[30]+4]<=REG[2];
      10'h212: data = 32'h8fc20008; // 00400848: LW, REG[2]<=RAM[REG[30]+8];
      10'h213: data = 32'h00000000; // 0040084c: SLL, REG[0]<=REG[0]<<0;
      10'h214: data = 32'h8c420000; // 00400850: LW, REG[2]<=RAM[REG[2]+0];
      10'h215: data = 32'h00000000; // 00400854: SLL, REG[0]<=REG[0]<<0;
      10'h216: data = 32'h2443ffd0; // 00400858: ADDIU, REG[3]<=REG[2]+65488(=0x0000ffd0);
      10'h217: data = 32'h8fc20004; // 0040085c: LW, REG[2]<=RAM[REG[30]+4];
      10'h218: data = 32'h00000000; // 00400860: SLL, REG[0]<=REG[0]<<0;
      10'h219: data = 32'h0043102b; // 00400864: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h21a: data = 32'h1440ffef; // 00400868: BNE, PC<=(REG[2] != REG[0])?PC+4+65519*4:PC+4;
      10'h21b: data = 32'h00000000; // 0040086c: SLL, REG[0]<=REG[0]<<0;
      10'h21c: data = 32'h8fc20008; // 00400870: LW, REG[2]<=RAM[REG[30]+8];
      10'h21d: data = 32'h00000000; // 00400874: SLL, REG[0]<=REG[0]<<0;
      10'h21e: data = 32'h24420004; // 00400878: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h21f: data = 32'hafc20008; // 0040087c: SW, RAM[REG[30]+8]<=REG[2];
      10'h220: data = 32'h8fc20008; // 00400880: LW, REG[2]<=RAM[REG[30]+8];
      10'h221: data = 32'h00000000; // 00400884: SLL, REG[0]<=REG[0]<<0;
      10'h222: data = 32'h8c430000; // 00400888: LW, REG[3]<=RAM[REG[2]+0];
      10'h223: data = 32'h8fc20000; // 0040088c: LW, REG[2]<=RAM[REG[30]+0];
      10'h224: data = 32'h00000000; // 00400890: SLL, REG[0]<=REG[0]<<0;
      10'h225: data = 32'h00621021; // 00400894: ADDU, REG[2]<=REG[3]+REG[2];
      10'h226: data = 32'h2442ffd0; // 00400898: ADDIU, REG[2]<=REG[2]+65488(=0x0000ffd0);
      10'h227: data = 32'hafc20000; // 0040089c: SW, RAM[REG[30]+0]<=REG[2];
      10'h228: data = 32'h8fc20000; // 004008a0: LW, REG[2]<=RAM[REG[30]+0];
      10'h229: data = 32'h03c0e821; // 004008a4: ADDU, REG[29]<=REG[30]+REG[0];
      10'h22a: data = 32'h8fbe0010; // 004008a8: LW, REG[30]<=RAM[REG[29]+16];
      10'h22b: data = 32'h27bd0018; // 004008ac: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h22c: data = 32'h03e00008; // 004008b0: JR, PC<=REG[31];
      10'h22d: data = 32'h00000000; // 004008b4: SLL, REG[0]<=REG[0]<<0;
      10'h22e: data = 32'h00000000; // 004008b8: SLL, REG[0]<=REG[0]<<0;
      10'h22f: data = 32'h00000000; // 004008bc: SLL, REG[0]<=REG[0]<<0;
    endcase
  end

  assign rom_data = data;
endmodule
