/*******************/
/* rom8x1024_sim.v */
/*******************/

//                  +----+
//  rom_addr[11:0]->|    |->rom_data[31:0]
//                  +----+

//
// ROM�ε��ҡ��������ߥ�졼������ѡ�
//

module rom8x1024_sim (rom_addr, rom_data);

  input   [11:0]  rom_addr;  // 12-bit ���ɥ쥹���ϥݡ���
  output  [31:0]  rom_data;  // 32-bit �ǡ������ϥݡ���

  reg     [31:0]  data;

  // Wire
  wire     [9:0]  word_addr; // 10-bit address, word

  assign word_addr = rom_addr[9:2];
   
  always @(word_addr) begin
    case (word_addr)
      10'h000: data = 32'he000001c; // 00400000: other type! opcode=56(10)
      10'h001: data = 32'h00000000; // 00400004: SLL, REG[0]<=REG[0]<<0;
      10'h002: data = 32'h00000000; // 00400008: SLL, REG[0]<=REG[0]<<0;
      10'h003: data = 32'h00000000; // 0040000c: SLL, REG[0]<=REG[0]<<0;
      10'h004: data = 32'h00000000; // 00400010: SLL, REG[0]<=REG[0]<<0;
      10'h005: data = 32'h00408800; // 00400014: SLL, REG[17]<=REG[0]<<0;
      10'h006: data = 32'h00000000; // 00400018: SLL, REG[0]<=REG[0]<<0;
      10'h007: data = 32'h00000000; // 0040001c: SLL, REG[0]<=REG[0]<<0;
      10'h008: data = 32'h27bdfee8; // 00400020: ADDIU, REG[29]<=REG[29]+65256(=0x0000fee8);
      10'h009: data = 32'hafbf0114; // 00400024: SW, RAM[REG[29]+276]<=REG[31];
      10'h00a: data = 32'hafbe0110; // 00400028: SW, RAM[REG[29]+272]<=REG[30];
      10'h00b: data = 32'h03a0f021; // 0040002c: ADDU, REG[30]<=REG[29]+REG[0];
      10'h00c: data = 32'h24020048; // 00400030: ADDIU, REG[2]<=REG[0]+72(=0x00000048);
      10'h00d: data = 32'hafc20010; // 00400034: SW, RAM[REG[30]+16]<=REG[2];
      10'h00e: data = 32'h24020045; // 00400038: ADDIU, REG[2]<=REG[0]+69(=0x00000045);
      10'h00f: data = 32'hafc20014; // 0040003c: SW, RAM[REG[30]+20]<=REG[2];
      10'h010: data = 32'h2402004c; // 00400040: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h011: data = 32'hafc20018; // 00400044: SW, RAM[REG[30]+24]<=REG[2];
      10'h012: data = 32'h2402004c; // 00400048: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h013: data = 32'hafc2001c; // 0040004c: SW, RAM[REG[30]+28]<=REG[2];
      10'h014: data = 32'h2402004f; // 00400050: ADDIU, REG[2]<=REG[0]+79(=0x0000004f);
      10'h015: data = 32'hafc20020; // 00400054: SW, RAM[REG[30]+32]<=REG[2];
      10'h016: data = 32'h24020021; // 00400058: ADDIU, REG[2]<=REG[0]+33(=0x00000021);
      10'h017: data = 32'hafc20024; // 0040005c: SW, RAM[REG[30]+36]<=REG[2];
      10'h018: data = 32'h24020021; // 00400060: ADDIU, REG[2]<=REG[0]+33(=0x00000021);
      10'h019: data = 32'hafc20028; // 00400064: SW, RAM[REG[30]+40]<=REG[2];
      10'h01a: data = 32'h2402000a; // 00400068: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h01b: data = 32'hafc2002c; // 0040006c: SW, RAM[REG[30]+44]<=REG[2];
      10'h01c: data = 32'hafc00030; // 00400070: SW, RAM[REG[30]+48]<=REG[0];
      10'h01d: data = 32'h27c20010; // 00400074: ADDIU, REG[2]<=REG[30]+16(=0x00000010);
      10'h01e: data = 32'h00402021; // 00400078: ADDU, REG[4]<=REG[2]+REG[0];
      10'h01f: data = 32'h0c100136; // 0040007c: JAL, PC<=0x00100136*4(=0x004004d8); REG[31]<=PC+4
      10'h020: data = 32'h00000000; // 00400080: SLL, REG[0]<=REG[0]<<0;
      10'h021: data = 32'h24020053; // 00400084: ADDIU, REG[2]<=REG[0]+83(=0x00000053);
      10'h022: data = 32'hafc20010; // 00400088: SW, RAM[REG[30]+16]<=REG[2];
      10'h023: data = 32'h24020054; // 0040008c: ADDIU, REG[2]<=REG[0]+84(=0x00000054);
      10'h024: data = 32'hafc20014; // 00400090: SW, RAM[REG[30]+20]<=REG[2];
      10'h025: data = 32'h24020052; // 00400094: ADDIU, REG[2]<=REG[0]+82(=0x00000052);
      10'h026: data = 32'hafc20018; // 00400098: SW, RAM[REG[30]+24]<=REG[2];
      10'h027: data = 32'h24020049; // 0040009c: ADDIU, REG[2]<=REG[0]+73(=0x00000049);
      10'h028: data = 32'hafc2001c; // 004000a0: SW, RAM[REG[30]+28]<=REG[2];
      10'h029: data = 32'h2402004e; // 004000a4: ADDIU, REG[2]<=REG[0]+78(=0x0000004e);
      10'h02a: data = 32'hafc20020; // 004000a8: SW, RAM[REG[30]+32]<=REG[2];
      10'h02b: data = 32'h24020047; // 004000ac: ADDIU, REG[2]<=REG[0]+71(=0x00000047);
      10'h02c: data = 32'hafc20024; // 004000b0: SW, RAM[REG[30]+36]<=REG[2];
      10'h02d: data = 32'h2402003d; // 004000b4: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h02e: data = 32'hafc20028; // 004000b8: SW, RAM[REG[30]+40]<=REG[2];
      10'h02f: data = 32'hafc0002c; // 004000bc: SW, RAM[REG[30]+44]<=REG[0];
      10'h030: data = 32'h27c20010; // 004000c0: ADDIU, REG[2]<=REG[30]+16(=0x00000010);
      10'h031: data = 32'h00402021; // 004000c4: ADDU, REG[4]<=REG[2]+REG[0];
      10'h032: data = 32'h0c100136; // 004000c8: JAL, PC<=0x00100136*4(=0x004004d8); REG[31]<=PC+4
      10'h033: data = 32'h00000000; // 004000cc: SLL, REG[0]<=REG[0]<<0;
      10'h034: data = 32'h27c20090; // 004000d0: ADDIU, REG[2]<=REG[30]+144(=0x00000090);
      10'h035: data = 32'h00402021; // 004000d4: ADDU, REG[4]<=REG[2]+REG[0];
      10'h036: data = 32'h0c100054; // 004000d8: JAL, PC<=0x00100054*4(=0x00400150); REG[31]<=PC+4
      10'h037: data = 32'h00000000; // 004000dc: SLL, REG[0]<=REG[0]<<0;
      10'h038: data = 32'h24020045; // 004000e0: ADDIU, REG[2]<=REG[0]+69(=0x00000045);
      10'h039: data = 32'hafc20010; // 004000e4: SW, RAM[REG[30]+16]<=REG[2];
      10'h03a: data = 32'h24020043; // 004000e8: ADDIU, REG[2]<=REG[0]+67(=0x00000043);
      10'h03b: data = 32'hafc20014; // 004000ec: SW, RAM[REG[30]+20]<=REG[2];
      10'h03c: data = 32'h24020048; // 004000f0: ADDIU, REG[2]<=REG[0]+72(=0x00000048);
      10'h03d: data = 32'hafc20018; // 004000f4: SW, RAM[REG[30]+24]<=REG[2];
      10'h03e: data = 32'h2402004f; // 004000f8: ADDIU, REG[2]<=REG[0]+79(=0x0000004f);
      10'h03f: data = 32'hafc2001c; // 004000fc: SW, RAM[REG[30]+28]<=REG[2];
      10'h040: data = 32'h24020020; // 00400100: ADDIU, REG[2]<=REG[0]+32(=0x00000020);
      10'h041: data = 32'hafc20020; // 00400104: SW, RAM[REG[30]+32]<=REG[2];
      10'h042: data = 32'hafc00024; // 00400108: SW, RAM[REG[30]+36]<=REG[0];
      10'h043: data = 32'h27c20010; // 0040010c: ADDIU, REG[2]<=REG[30]+16(=0x00000010);
      10'h044: data = 32'h00402021; // 00400110: ADDU, REG[4]<=REG[2]+REG[0];
      10'h045: data = 32'h0c100136; // 00400114: JAL, PC<=0x00100136*4(=0x004004d8); REG[31]<=PC+4
      10'h046: data = 32'h00000000; // 00400118: SLL, REG[0]<=REG[0]<<0;
      10'h047: data = 32'h27c20090; // 0040011c: ADDIU, REG[2]<=REG[30]+144(=0x00000090);
      10'h048: data = 32'h00402021; // 00400120: ADDU, REG[4]<=REG[2]+REG[0];
      10'h049: data = 32'h0c100136; // 00400124: JAL, PC<=0x00100136*4(=0x004004d8); REG[31]<=PC+4
      10'h04a: data = 32'h00000000; // 00400128: SLL, REG[0]<=REG[0]<<0;
      10'h04b: data = 32'h2402000a; // 0040012c: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h04c: data = 32'hafc20010; // 00400130: SW, RAM[REG[30]+16]<=REG[2];
      10'h04d: data = 32'hafc00014; // 00400134: SW, RAM[REG[30]+20]<=REG[0];
      10'h04e: data = 32'h27c20010; // 00400138: ADDIU, REG[2]<=REG[30]+16(=0x00000010);
      10'h04f: data = 32'h00402021; // 0040013c: ADDU, REG[4]<=REG[2]+REG[0];
      10'h050: data = 32'h0c100136; // 00400140: JAL, PC<=0x00100136*4(=0x004004d8); REG[31]<=PC+4
      10'h051: data = 32'h00000000; // 00400144: SLL, REG[0]<=REG[0]<<0;
      10'h052: data = 32'h08100021; // 00400148: J, PC<=0x00100021*4(=0x00400084);
      10'h053: data = 32'h00000000; // 0040014c: SLL, REG[0]<=REG[0]<<0;
      10'h054: data = 32'h27bdfff8; // 00400150: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h055: data = 32'hafbe0000; // 00400154: SW, RAM[REG[29]+0]<=REG[30];
      10'h056: data = 32'h03a0f021; // 00400158: ADDU, REG[30]<=REG[29]+REG[0];
      10'h057: data = 32'hafc40008; // 0040015c: SW, RAM[REG[30]+8]<=REG[4];
      10'h058: data = 32'h24020308; // 00400160: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h059: data = 32'hac400000; // 00400164: SW, RAM[REG[2]+0]<=REG[0];
      10'h05a: data = 32'h2403030c; // 00400168: ADDIU, REG[3]<=REG[0]+780(=0x0000030c);
      10'h05b: data = 32'h24020001; // 0040016c: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h05c: data = 32'hac620000; // 00400170: SW, RAM[REG[3]+0]<=REG[2];
      10'h05d: data = 32'h24030308; // 00400174: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h05e: data = 32'h24020001; // 00400178: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h05f: data = 32'hac620000; // 0040017c: SW, RAM[REG[3]+0]<=REG[2];
      10'h060: data = 32'h24020308; // 00400180: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h061: data = 32'hac400000; // 00400184: SW, RAM[REG[2]+0]<=REG[0];
      10'h062: data = 32'h24030308; // 00400188: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h063: data = 32'h24020001; // 0040018c: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h064: data = 32'hac620000; // 00400190: SW, RAM[REG[3]+0]<=REG[2];
      10'h065: data = 32'h0810006c; // 00400194: J, PC<=0x0010006c*4(=0x004001b0);
      10'h066: data = 32'h00000000; // 00400198: SLL, REG[0]<=REG[0]<<0;
      10'h067: data = 32'h24020308; // 0040019c: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h068: data = 32'hac400000; // 004001a0: SW, RAM[REG[2]+0]<=REG[0];
      10'h069: data = 32'h24030308; // 004001a4: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h06a: data = 32'h24020001; // 004001a8: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h06b: data = 32'hac620000; // 004001ac: SW, RAM[REG[3]+0]<=REG[2];
      10'h06c: data = 32'h24020310; // 004001b0: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h06d: data = 32'h8c430000; // 004001b4: LW, REG[3]<=RAM[REG[2]+0];
      10'h06e: data = 32'h2402ffff; // 004001b8: ADDIU, REG[2]<=REG[0]+65535(=0x0000ffff);
      10'h06f: data = 32'h1062fff7; // 004001bc: BEQ, PC<=(REG[3] == REG[2])?PC+4+65527*4:PC+4;
      10'h070: data = 32'h00000000; // 004001c0: SLL, REG[0]<=REG[0]<<0;
      10'h071: data = 32'h0810011a; // 004001c4: J, PC<=0x0010011a*4(=0x00400468);
      10'h072: data = 32'h00000000; // 004001c8: SLL, REG[0]<=REG[0]<<0;
      10'h073: data = 32'h8fc20008; // 004001cc: LW, REG[2]<=RAM[REG[30]+8];
      10'h074: data = 32'h00000000; // 004001d0: SLL, REG[0]<=REG[0]<<0;
      10'h075: data = 32'h8c420000; // 004001d4: LW, REG[2]<=RAM[REG[2]+0];
      10'h076: data = 32'h00000000; // 004001d8: SLL, REG[0]<=REG[0]<<0;
      10'h077: data = 32'h10400012; // 004001dc: BEQ, PC<=(REG[2] == REG[0])?PC+4+18*4:PC+4;
      10'h078: data = 32'h00000000; // 004001e0: SLL, REG[0]<=REG[0]<<0;
      10'h079: data = 32'h8fc20008; // 004001e4: LW, REG[2]<=RAM[REG[30]+8];
      10'h07a: data = 32'h00000000; // 004001e8: SLL, REG[0]<=REG[0]<<0;
      10'h07b: data = 32'h8c420000; // 004001ec: LW, REG[2]<=RAM[REG[2]+0];
      10'h07c: data = 32'h00000000; // 004001f0: SLL, REG[0]<=REG[0]<<0;
      10'h07d: data = 32'h2c42001b; // 004001f4: SLTIU, REG[2]<=(REG[2]<27(=0x0000001b))?1:0;
      10'h07e: data = 32'h1040000b; // 004001f8: BEQ, PC<=(REG[2] == REG[0])?PC+4+11*4:PC+4;
      10'h07f: data = 32'h00000000; // 004001fc: SLL, REG[0]<=REG[0]<<0;
      10'h080: data = 32'h8fc20008; // 00400200: LW, REG[2]<=RAM[REG[30]+8];
      10'h081: data = 32'h00000000; // 00400204: SLL, REG[0]<=REG[0]<<0;
      10'h082: data = 32'h8c420000; // 00400208: LW, REG[2]<=RAM[REG[2]+0];
      10'h083: data = 32'h00000000; // 0040020c: SLL, REG[0]<=REG[0]<<0;
      10'h084: data = 32'h24430040; // 00400210: ADDIU, REG[3]<=REG[2]+64(=0x00000040);
      10'h085: data = 32'h8fc20008; // 00400214: LW, REG[2]<=RAM[REG[30]+8];
      10'h086: data = 32'h00000000; // 00400218: SLL, REG[0]<=REG[0]<<0;
      10'h087: data = 32'hac430000; // 0040021c: SW, RAM[REG[2]+0]<=REG[3];
      10'h088: data = 32'h08100111; // 00400220: J, PC<=0x00100111*4(=0x00400444);
      10'h089: data = 32'h00000000; // 00400224: SLL, REG[0]<=REG[0]<<0;
      10'h08a: data = 32'h8fc20008; // 00400228: LW, REG[2]<=RAM[REG[30]+8];
      10'h08b: data = 32'h00000000; // 0040022c: SLL, REG[0]<=REG[0]<<0;
      10'h08c: data = 32'h8c420000; // 00400230: LW, REG[2]<=RAM[REG[2]+0];
      10'h08d: data = 32'h00000000; // 00400234: SLL, REG[0]<=REG[0]<<0;
      10'h08e: data = 32'h2c420030; // 00400238: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h08f: data = 32'h14400010; // 0040023c: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h090: data = 32'h00000000; // 00400240: SLL, REG[0]<=REG[0]<<0;
      10'h091: data = 32'h8fc20008; // 00400244: LW, REG[2]<=RAM[REG[30]+8];
      10'h092: data = 32'h00000000; // 00400248: SLL, REG[0]<=REG[0]<<0;
      10'h093: data = 32'h8c420000; // 0040024c: LW, REG[2]<=RAM[REG[2]+0];
      10'h094: data = 32'h00000000; // 00400250: SLL, REG[0]<=REG[0]<<0;
      10'h095: data = 32'h2c42003a; // 00400254: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h096: data = 32'h10400009; // 00400258: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h097: data = 32'h00000000; // 0040025c: SLL, REG[0]<=REG[0]<<0;
      10'h098: data = 32'h8fc20008; // 00400260: LW, REG[2]<=RAM[REG[30]+8];
      10'h099: data = 32'h00000000; // 00400264: SLL, REG[0]<=REG[0]<<0;
      10'h09a: data = 32'h8c430000; // 00400268: LW, REG[3]<=RAM[REG[2]+0];
      10'h09b: data = 32'h8fc20008; // 0040026c: LW, REG[2]<=RAM[REG[30]+8];
      10'h09c: data = 32'h00000000; // 00400270: SLL, REG[0]<=REG[0]<<0;
      10'h09d: data = 32'hac430000; // 00400274: SW, RAM[REG[2]+0]<=REG[3];
      10'h09e: data = 32'h08100111; // 00400278: J, PC<=0x00100111*4(=0x00400444);
      10'h09f: data = 32'h00000000; // 0040027c: SLL, REG[0]<=REG[0]<<0;
      10'h0a0: data = 32'h8fc20008; // 00400280: LW, REG[2]<=RAM[REG[30]+8];
      10'h0a1: data = 32'h00000000; // 00400284: SLL, REG[0]<=REG[0]<<0;
      10'h0a2: data = 32'h8c420000; // 00400288: LW, REG[2]<=RAM[REG[2]+0];
      10'h0a3: data = 32'h00000000; // 0040028c: SLL, REG[0]<=REG[0]<<0;
      10'h0a4: data = 32'h14400006; // 00400290: BNE, PC<=(REG[2] != REG[0])?PC+4+6*4:PC+4;
      10'h0a5: data = 32'h00000000; // 00400294: SLL, REG[0]<=REG[0]<<0;
      10'h0a6: data = 32'h8fc30008; // 00400298: LW, REG[3]<=RAM[REG[30]+8];
      10'h0a7: data = 32'h24020040; // 0040029c: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h0a8: data = 32'hac620000; // 004002a0: SW, RAM[REG[3]+0]<=REG[2];
      10'h0a9: data = 32'h08100111; // 004002a4: J, PC<=0x00100111*4(=0x00400444);
      10'h0aa: data = 32'h00000000; // 004002a8: SLL, REG[0]<=REG[0]<<0;
      10'h0ab: data = 32'h8fc20008; // 004002ac: LW, REG[2]<=RAM[REG[30]+8];
      10'h0ac: data = 32'h00000000; // 004002b0: SLL, REG[0]<=REG[0]<<0;
      10'h0ad: data = 32'h8c430000; // 004002b4: LW, REG[3]<=RAM[REG[2]+0];
      10'h0ae: data = 32'h2402001b; // 004002b8: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h0af: data = 32'h14620006; // 004002bc: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0b0: data = 32'h00000000; // 004002c0: SLL, REG[0]<=REG[0]<<0;
      10'h0b1: data = 32'h8fc30008; // 004002c4: LW, REG[3]<=RAM[REG[30]+8];
      10'h0b2: data = 32'h2402005b; // 004002c8: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h0b3: data = 32'hac620000; // 004002cc: SW, RAM[REG[3]+0]<=REG[2];
      10'h0b4: data = 32'h08100111; // 004002d0: J, PC<=0x00100111*4(=0x00400444);
      10'h0b5: data = 32'h00000000; // 004002d4: SLL, REG[0]<=REG[0]<<0;
      10'h0b6: data = 32'h8fc20008; // 004002d8: LW, REG[2]<=RAM[REG[30]+8];
      10'h0b7: data = 32'h00000000; // 004002dc: SLL, REG[0]<=REG[0]<<0;
      10'h0b8: data = 32'h8c430000; // 004002e0: LW, REG[3]<=RAM[REG[2]+0];
      10'h0b9: data = 32'h2402001d; // 004002e4: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h0ba: data = 32'h14620006; // 004002e8: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0bb: data = 32'h00000000; // 004002ec: SLL, REG[0]<=REG[0]<<0;
      10'h0bc: data = 32'h8fc30008; // 004002f0: LW, REG[3]<=RAM[REG[30]+8];
      10'h0bd: data = 32'h2402005d; // 004002f4: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h0be: data = 32'hac620000; // 004002f8: SW, RAM[REG[3]+0]<=REG[2];
      10'h0bf: data = 32'h08100111; // 004002fc: J, PC<=0x00100111*4(=0x00400444);
      10'h0c0: data = 32'h00000000; // 00400300: SLL, REG[0]<=REG[0]<<0;
      10'h0c1: data = 32'h8fc20008; // 00400304: LW, REG[2]<=RAM[REG[30]+8];
      10'h0c2: data = 32'h00000000; // 00400308: SLL, REG[0]<=REG[0]<<0;
      10'h0c3: data = 32'h8c420000; // 0040030c: LW, REG[2]<=RAM[REG[2]+0];
      10'h0c4: data = 32'h00000000; // 00400310: SLL, REG[0]<=REG[0]<<0;
      10'h0c5: data = 32'h2c420020; // 00400314: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h0c6: data = 32'h14400010; // 00400318: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h0c7: data = 32'h00000000; // 0040031c: SLL, REG[0]<=REG[0]<<0;
      10'h0c8: data = 32'h8fc20008; // 00400320: LW, REG[2]<=RAM[REG[30]+8];
      10'h0c9: data = 32'h00000000; // 00400324: SLL, REG[0]<=REG[0]<<0;
      10'h0ca: data = 32'h8c420000; // 00400328: LW, REG[2]<=RAM[REG[2]+0];
      10'h0cb: data = 32'h00000000; // 0040032c: SLL, REG[0]<=REG[0]<<0;
      10'h0cc: data = 32'h2c420030; // 00400330: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h0cd: data = 32'h10400009; // 00400334: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h0ce: data = 32'h00000000; // 00400338: SLL, REG[0]<=REG[0]<<0;
      10'h0cf: data = 32'h8fc20008; // 0040033c: LW, REG[2]<=RAM[REG[30]+8];
      10'h0d0: data = 32'h00000000; // 00400340: SLL, REG[0]<=REG[0]<<0;
      10'h0d1: data = 32'h8c430000; // 00400344: LW, REG[3]<=RAM[REG[2]+0];
      10'h0d2: data = 32'h8fc20008; // 00400348: LW, REG[2]<=RAM[REG[30]+8];
      10'h0d3: data = 32'h00000000; // 0040034c: SLL, REG[0]<=REG[0]<<0;
      10'h0d4: data = 32'hac430000; // 00400350: SW, RAM[REG[2]+0]<=REG[3];
      10'h0d5: data = 32'h08100111; // 00400354: J, PC<=0x00100111*4(=0x00400444);
      10'h0d6: data = 32'h00000000; // 00400358: SLL, REG[0]<=REG[0]<<0;
      10'h0d7: data = 32'h8fc20008; // 0040035c: LW, REG[2]<=RAM[REG[30]+8];
      10'h0d8: data = 32'h00000000; // 00400360: SLL, REG[0]<=REG[0]<<0;
      10'h0d9: data = 32'h8c430000; // 00400364: LW, REG[3]<=RAM[REG[2]+0];
      10'h0da: data = 32'h2402003a; // 00400368: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h0db: data = 32'h14620006; // 0040036c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0dc: data = 32'h00000000; // 00400370: SLL, REG[0]<=REG[0]<<0;
      10'h0dd: data = 32'h8fc30008; // 00400374: LW, REG[3]<=RAM[REG[30]+8];
      10'h0de: data = 32'h2402003f; // 00400378: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h0df: data = 32'hac620000; // 0040037c: SW, RAM[REG[3]+0]<=REG[2];
      10'h0e0: data = 32'h08100111; // 00400380: J, PC<=0x00100111*4(=0x00400444);
      10'h0e1: data = 32'h00000000; // 00400384: SLL, REG[0]<=REG[0]<<0;
      10'h0e2: data = 32'h8fc20008; // 00400388: LW, REG[2]<=RAM[REG[30]+8];
      10'h0e3: data = 32'h00000000; // 0040038c: SLL, REG[0]<=REG[0]<<0;
      10'h0e4: data = 32'h8c430000; // 00400390: LW, REG[3]<=RAM[REG[2]+0];
      10'h0e5: data = 32'h2402003b; // 00400394: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h0e6: data = 32'h14620006; // 00400398: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0e7: data = 32'h00000000; // 0040039c: SLL, REG[0]<=REG[0]<<0;
      10'h0e8: data = 32'h8fc30008; // 004003a0: LW, REG[3]<=RAM[REG[30]+8];
      10'h0e9: data = 32'h2402003d; // 004003a4: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h0ea: data = 32'hac620000; // 004003a8: SW, RAM[REG[3]+0]<=REG[2];
      10'h0eb: data = 32'h08100111; // 004003ac: J, PC<=0x00100111*4(=0x00400444);
      10'h0ec: data = 32'h00000000; // 004003b0: SLL, REG[0]<=REG[0]<<0;
      10'h0ed: data = 32'h8fc20008; // 004003b4: LW, REG[2]<=RAM[REG[30]+8];
      10'h0ee: data = 32'h00000000; // 004003b8: SLL, REG[0]<=REG[0]<<0;
      10'h0ef: data = 32'h8c430000; // 004003bc: LW, REG[3]<=RAM[REG[2]+0];
      10'h0f0: data = 32'h2402003c; // 004003c0: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h0f1: data = 32'h14620006; // 004003c4: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0f2: data = 32'h00000000; // 004003c8: SLL, REG[0]<=REG[0]<<0;
      10'h0f3: data = 32'h8fc30008; // 004003cc: LW, REG[3]<=RAM[REG[30]+8];
      10'h0f4: data = 32'h2402003b; // 004003d0: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h0f5: data = 32'hac620000; // 004003d4: SW, RAM[REG[3]+0]<=REG[2];
      10'h0f6: data = 32'h08100111; // 004003d8: J, PC<=0x00100111*4(=0x00400444);
      10'h0f7: data = 32'h00000000; // 004003dc: SLL, REG[0]<=REG[0]<<0;
      10'h0f8: data = 32'h8fc20008; // 004003e0: LW, REG[2]<=RAM[REG[30]+8];
      10'h0f9: data = 32'h00000000; // 004003e4: SLL, REG[0]<=REG[0]<<0;
      10'h0fa: data = 32'h8c430000; // 004003e8: LW, REG[3]<=RAM[REG[2]+0];
      10'h0fb: data = 32'h2402003d; // 004003ec: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h0fc: data = 32'h14620006; // 004003f0: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0fd: data = 32'h00000000; // 004003f4: SLL, REG[0]<=REG[0]<<0;
      10'h0fe: data = 32'h8fc30008; // 004003f8: LW, REG[3]<=RAM[REG[30]+8];
      10'h0ff: data = 32'h2402003a; // 004003fc: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h100: data = 32'hac620000; // 00400400: SW, RAM[REG[3]+0]<=REG[2];
      10'h101: data = 32'h08100111; // 00400404: J, PC<=0x00100111*4(=0x00400444);
      10'h102: data = 32'h00000000; // 00400408: SLL, REG[0]<=REG[0]<<0;
      10'h103: data = 32'h8fc20008; // 0040040c: LW, REG[2]<=RAM[REG[30]+8];
      10'h104: data = 32'h00000000; // 00400410: SLL, REG[0]<=REG[0]<<0;
      10'h105: data = 32'h8c430000; // 00400414: LW, REG[3]<=RAM[REG[2]+0];
      10'h106: data = 32'h2402003e; // 00400418: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h107: data = 32'h14620006; // 0040041c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h108: data = 32'h00000000; // 00400420: SLL, REG[0]<=REG[0]<<0;
      10'h109: data = 32'h8fc30008; // 00400424: LW, REG[3]<=RAM[REG[30]+8];
      10'h10a: data = 32'h2402000a; // 00400428: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h10b: data = 32'hac620000; // 0040042c: SW, RAM[REG[3]+0]<=REG[2];
      10'h10c: data = 32'h08100111; // 00400430: J, PC<=0x00100111*4(=0x00400444);
      10'h10d: data = 32'h00000000; // 00400434: SLL, REG[0]<=REG[0]<<0;
      10'h10e: data = 32'h8fc30008; // 00400438: LW, REG[3]<=RAM[REG[30]+8];
      10'h10f: data = 32'h24020040; // 0040043c: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h110: data = 32'hac620000; // 00400440: SW, RAM[REG[3]+0]<=REG[2];
      10'h111: data = 32'h24020308; // 00400444: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h112: data = 32'hac400000; // 00400448: SW, RAM[REG[2]+0]<=REG[0];
      10'h113: data = 32'h24030308; // 0040044c: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h114: data = 32'h24020001; // 00400450: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h115: data = 32'hac620000; // 00400454: SW, RAM[REG[3]+0]<=REG[2];
      10'h116: data = 32'h8fc20008; // 00400458: LW, REG[2]<=RAM[REG[30]+8];
      10'h117: data = 32'h00000000; // 0040045c: SLL, REG[0]<=REG[0]<<0;
      10'h118: data = 32'h24420004; // 00400460: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h119: data = 32'hafc20008; // 00400464: SW, RAM[REG[30]+8]<=REG[2];
      10'h11a: data = 32'h24020310; // 00400468: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h11b: data = 32'h8c430000; // 0040046c: LW, REG[3]<=RAM[REG[2]+0];
      10'h11c: data = 32'h8fc20008; // 00400470: LW, REG[2]<=RAM[REG[30]+8];
      10'h11d: data = 32'h00000000; // 00400474: SLL, REG[0]<=REG[0]<<0;
      10'h11e: data = 32'hac430000; // 00400478: SW, RAM[REG[2]+0]<=REG[3];
      10'h11f: data = 32'h8fc20008; // 0040047c: LW, REG[2]<=RAM[REG[30]+8];
      10'h120: data = 32'h00000000; // 00400480: SLL, REG[0]<=REG[0]<<0;
      10'h121: data = 32'h8c430000; // 00400484: LW, REG[3]<=RAM[REG[2]+0];
      10'h122: data = 32'h2402003e; // 00400488: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h123: data = 32'h1462ff4f; // 0040048c: BNE, PC<=(REG[3] != REG[2])?PC+4+65359*4:PC+4;
      10'h124: data = 32'h00000000; // 00400490: SLL, REG[0]<=REG[0]<<0;
      10'h125: data = 32'h8fc20008; // 00400494: LW, REG[2]<=RAM[REG[30]+8];
      10'h126: data = 32'h00000000; // 00400498: SLL, REG[0]<=REG[0]<<0;
      10'h127: data = 32'hac400000; // 0040049c: SW, RAM[REG[2]+0]<=REG[0];
      10'h128: data = 32'h24020308; // 004004a0: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h129: data = 32'hac400000; // 004004a4: SW, RAM[REG[2]+0]<=REG[0];
      10'h12a: data = 32'h2402030c; // 004004a8: ADDIU, REG[2]<=REG[0]+780(=0x0000030c);
      10'h12b: data = 32'hac400000; // 004004ac: SW, RAM[REG[2]+0]<=REG[0];
      10'h12c: data = 32'h24030308; // 004004b0: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h12d: data = 32'h24020001; // 004004b4: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h12e: data = 32'hac620000; // 004004b8: SW, RAM[REG[3]+0]<=REG[2];
      10'h12f: data = 32'h24020308; // 004004bc: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h130: data = 32'hac400000; // 004004c0: SW, RAM[REG[2]+0]<=REG[0];
      10'h131: data = 32'h03c0e821; // 004004c4: ADDU, REG[29]<=REG[30]+REG[0];
      10'h132: data = 32'h8fbe0000; // 004004c8: LW, REG[30]<=RAM[REG[29]+0];
      10'h133: data = 32'h27bd0008; // 004004cc: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h134: data = 32'h03e00008; // 004004d0: JR, PC<=REG[31];
      10'h135: data = 32'h00000000; // 004004d4: SLL, REG[0]<=REG[0]<<0;
      10'h136: data = 32'h27bdfff8; // 004004d8: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h137: data = 32'hafbe0000; // 004004dc: SW, RAM[REG[29]+0]<=REG[30];
      10'h138: data = 32'h03a0f021; // 004004e0: ADDU, REG[30]<=REG[29]+REG[0];
      10'h139: data = 32'hafc40008; // 004004e4: SW, RAM[REG[30]+8]<=REG[4];
      10'h13a: data = 32'h081001f8; // 004004e8: J, PC<=0x001001f8*4(=0x004007e0);
      10'h13b: data = 32'h00000000; // 004004ec: SLL, REG[0]<=REG[0]<<0;
      10'h13c: data = 32'h24020300; // 004004f0: ADDIU, REG[2]<=REG[0]+768(=0x00000300);
      10'h13d: data = 32'hac400000; // 004004f4: SW, RAM[REG[2]+0]<=REG[0];
      10'h13e: data = 32'h8fc20008; // 004004f8: LW, REG[2]<=RAM[REG[30]+8];
      10'h13f: data = 32'h00000000; // 004004fc: SLL, REG[0]<=REG[0]<<0;
      10'h140: data = 32'h8c420000; // 00400500: LW, REG[2]<=RAM[REG[2]+0];
      10'h141: data = 32'h00000000; // 00400504: SLL, REG[0]<=REG[0]<<0;
      10'h142: data = 32'h2c420041; // 00400508: SLTIU, REG[2]<=(REG[2]<65(=0x00000041))?1:0;
      10'h143: data = 32'h14400011; // 0040050c: BNE, PC<=(REG[2] != REG[0])?PC+4+17*4:PC+4;
      10'h144: data = 32'h00000000; // 00400510: SLL, REG[0]<=REG[0]<<0;
      10'h145: data = 32'h8fc20008; // 00400514: LW, REG[2]<=RAM[REG[30]+8];
      10'h146: data = 32'h00000000; // 00400518: SLL, REG[0]<=REG[0]<<0;
      10'h147: data = 32'h8c420000; // 0040051c: LW, REG[2]<=RAM[REG[2]+0];
      10'h148: data = 32'h00000000; // 00400520: SLL, REG[0]<=REG[0]<<0;
      10'h149: data = 32'h2c42005b; // 00400524: SLTIU, REG[2]<=(REG[2]<91(=0x0000005b))?1:0;
      10'h14a: data = 32'h1040000a; // 00400528: BEQ, PC<=(REG[2] == REG[0])?PC+4+10*4:PC+4;
      10'h14b: data = 32'h00000000; // 0040052c: SLL, REG[0]<=REG[0]<<0;
      10'h14c: data = 32'h24030304; // 00400530: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h14d: data = 32'h8fc20008; // 00400534: LW, REG[2]<=RAM[REG[30]+8];
      10'h14e: data = 32'h00000000; // 00400538: SLL, REG[0]<=REG[0]<<0;
      10'h14f: data = 32'h8c420000; // 0040053c: LW, REG[2]<=RAM[REG[2]+0];
      10'h150: data = 32'h00000000; // 00400540: SLL, REG[0]<=REG[0]<<0;
      10'h151: data = 32'h2442ffc0; // 00400544: ADDIU, REG[2]<=REG[2]+65472(=0x0000ffc0);
      10'h152: data = 32'hac620000; // 00400548: SW, RAM[REG[3]+0]<=REG[2];
      10'h153: data = 32'h081001f1; // 0040054c: J, PC<=0x001001f1*4(=0x004007c4);
      10'h154: data = 32'h00000000; // 00400550: SLL, REG[0]<=REG[0]<<0;
      10'h155: data = 32'h8fc20008; // 00400554: LW, REG[2]<=RAM[REG[30]+8];
      10'h156: data = 32'h00000000; // 00400558: SLL, REG[0]<=REG[0]<<0;
      10'h157: data = 32'h8c420000; // 0040055c: LW, REG[2]<=RAM[REG[2]+0];
      10'h158: data = 32'h00000000; // 00400560: SLL, REG[0]<=REG[0]<<0;
      10'h159: data = 32'h2c420061; // 00400564: SLTIU, REG[2]<=(REG[2]<97(=0x00000061))?1:0;
      10'h15a: data = 32'h14400011; // 00400568: BNE, PC<=(REG[2] != REG[0])?PC+4+17*4:PC+4;
      10'h15b: data = 32'h00000000; // 0040056c: SLL, REG[0]<=REG[0]<<0;
      10'h15c: data = 32'h8fc20008; // 00400570: LW, REG[2]<=RAM[REG[30]+8];
      10'h15d: data = 32'h00000000; // 00400574: SLL, REG[0]<=REG[0]<<0;
      10'h15e: data = 32'h8c420000; // 00400578: LW, REG[2]<=RAM[REG[2]+0];
      10'h15f: data = 32'h00000000; // 0040057c: SLL, REG[0]<=REG[0]<<0;
      10'h160: data = 32'h2c42007b; // 00400580: SLTIU, REG[2]<=(REG[2]<123(=0x0000007b))?1:0;
      10'h161: data = 32'h1040000a; // 00400584: BEQ, PC<=(REG[2] == REG[0])?PC+4+10*4:PC+4;
      10'h162: data = 32'h00000000; // 00400588: SLL, REG[0]<=REG[0]<<0;
      10'h163: data = 32'h24030304; // 0040058c: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h164: data = 32'h8fc20008; // 00400590: LW, REG[2]<=RAM[REG[30]+8];
      10'h165: data = 32'h00000000; // 00400594: SLL, REG[0]<=REG[0]<<0;
      10'h166: data = 32'h8c420000; // 00400598: LW, REG[2]<=RAM[REG[2]+0];
      10'h167: data = 32'h00000000; // 0040059c: SLL, REG[0]<=REG[0]<<0;
      10'h168: data = 32'h2442ffa0; // 004005a0: ADDIU, REG[2]<=REG[2]+65440(=0x0000ffa0);
      10'h169: data = 32'hac620000; // 004005a4: SW, RAM[REG[3]+0]<=REG[2];
      10'h16a: data = 32'h081001f1; // 004005a8: J, PC<=0x001001f1*4(=0x004007c4);
      10'h16b: data = 32'h00000000; // 004005ac: SLL, REG[0]<=REG[0]<<0;
      10'h16c: data = 32'h8fc20008; // 004005b0: LW, REG[2]<=RAM[REG[30]+8];
      10'h16d: data = 32'h00000000; // 004005b4: SLL, REG[0]<=REG[0]<<0;
      10'h16e: data = 32'h8c420000; // 004005b8: LW, REG[2]<=RAM[REG[2]+0];
      10'h16f: data = 32'h00000000; // 004005bc: SLL, REG[0]<=REG[0]<<0;
      10'h170: data = 32'h2c420030; // 004005c0: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h171: data = 32'h14400010; // 004005c4: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h172: data = 32'h00000000; // 004005c8: SLL, REG[0]<=REG[0]<<0;
      10'h173: data = 32'h8fc20008; // 004005cc: LW, REG[2]<=RAM[REG[30]+8];
      10'h174: data = 32'h00000000; // 004005d0: SLL, REG[0]<=REG[0]<<0;
      10'h175: data = 32'h8c420000; // 004005d4: LW, REG[2]<=RAM[REG[2]+0];
      10'h176: data = 32'h00000000; // 004005d8: SLL, REG[0]<=REG[0]<<0;
      10'h177: data = 32'h2c42003a; // 004005dc: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h178: data = 32'h10400009; // 004005e0: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h179: data = 32'h00000000; // 004005e4: SLL, REG[0]<=REG[0]<<0;
      10'h17a: data = 32'h24020304; // 004005e8: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h17b: data = 32'h8fc30008; // 004005ec: LW, REG[3]<=RAM[REG[30]+8];
      10'h17c: data = 32'h00000000; // 004005f0: SLL, REG[0]<=REG[0]<<0;
      10'h17d: data = 32'h8c630000; // 004005f4: LW, REG[3]<=RAM[REG[3]+0];
      10'h17e: data = 32'h00000000; // 004005f8: SLL, REG[0]<=REG[0]<<0;
      10'h17f: data = 32'hac430000; // 004005fc: SW, RAM[REG[2]+0]<=REG[3];
      10'h180: data = 32'h081001f1; // 00400600: J, PC<=0x001001f1*4(=0x004007c4);
      10'h181: data = 32'h00000000; // 00400604: SLL, REG[0]<=REG[0]<<0;
      10'h182: data = 32'h8fc20008; // 00400608: LW, REG[2]<=RAM[REG[30]+8];
      10'h183: data = 32'h00000000; // 0040060c: SLL, REG[0]<=REG[0]<<0;
      10'h184: data = 32'h8c430000; // 00400610: LW, REG[3]<=RAM[REG[2]+0];
      10'h185: data = 32'h24020040; // 00400614: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h186: data = 32'h14620005; // 00400618: BNE, PC<=(REG[3] != REG[2])?PC+4+5*4:PC+4;
      10'h187: data = 32'h00000000; // 0040061c: SLL, REG[0]<=REG[0]<<0;
      10'h188: data = 32'h24020304; // 00400620: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h189: data = 32'hac400000; // 00400624: SW, RAM[REG[2]+0]<=REG[0];
      10'h18a: data = 32'h081001f1; // 00400628: J, PC<=0x001001f1*4(=0x004007c4);
      10'h18b: data = 32'h00000000; // 0040062c: SLL, REG[0]<=REG[0]<<0;
      10'h18c: data = 32'h8fc20008; // 00400630: LW, REG[2]<=RAM[REG[30]+8];
      10'h18d: data = 32'h00000000; // 00400634: SLL, REG[0]<=REG[0]<<0;
      10'h18e: data = 32'h8c430000; // 00400638: LW, REG[3]<=RAM[REG[2]+0];
      10'h18f: data = 32'h2402005b; // 0040063c: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h190: data = 32'h14620006; // 00400640: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h191: data = 32'h00000000; // 00400644: SLL, REG[0]<=REG[0]<<0;
      10'h192: data = 32'h24030304; // 00400648: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h193: data = 32'h2402001b; // 0040064c: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h194: data = 32'hac620000; // 00400650: SW, RAM[REG[3]+0]<=REG[2];
      10'h195: data = 32'h081001f1; // 00400654: J, PC<=0x001001f1*4(=0x004007c4);
      10'h196: data = 32'h00000000; // 00400658: SLL, REG[0]<=REG[0]<<0;
      10'h197: data = 32'h8fc20008; // 0040065c: LW, REG[2]<=RAM[REG[30]+8];
      10'h198: data = 32'h00000000; // 00400660: SLL, REG[0]<=REG[0]<<0;
      10'h199: data = 32'h8c430000; // 00400664: LW, REG[3]<=RAM[REG[2]+0];
      10'h19a: data = 32'h2402005d; // 00400668: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h19b: data = 32'h14620006; // 0040066c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h19c: data = 32'h00000000; // 00400670: SLL, REG[0]<=REG[0]<<0;
      10'h19d: data = 32'h24030304; // 00400674: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h19e: data = 32'h2402001d; // 00400678: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h19f: data = 32'hac620000; // 0040067c: SW, RAM[REG[3]+0]<=REG[2];
      10'h1a0: data = 32'h081001f1; // 00400680: J, PC<=0x001001f1*4(=0x004007c4);
      10'h1a1: data = 32'h00000000; // 00400684: SLL, REG[0]<=REG[0]<<0;
      10'h1a2: data = 32'h8fc20008; // 00400688: LW, REG[2]<=RAM[REG[30]+8];
      10'h1a3: data = 32'h00000000; // 0040068c: SLL, REG[0]<=REG[0]<<0;
      10'h1a4: data = 32'h8c420000; // 00400690: LW, REG[2]<=RAM[REG[2]+0];
      10'h1a5: data = 32'h00000000; // 00400694: SLL, REG[0]<=REG[0]<<0;
      10'h1a6: data = 32'h2c420020; // 00400698: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h1a7: data = 32'h14400010; // 0040069c: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h1a8: data = 32'h00000000; // 004006a0: SLL, REG[0]<=REG[0]<<0;
      10'h1a9: data = 32'h8fc20008; // 004006a4: LW, REG[2]<=RAM[REG[30]+8];
      10'h1aa: data = 32'h00000000; // 004006a8: SLL, REG[0]<=REG[0]<<0;
      10'h1ab: data = 32'h8c420000; // 004006ac: LW, REG[2]<=RAM[REG[2]+0];
      10'h1ac: data = 32'h00000000; // 004006b0: SLL, REG[0]<=REG[0]<<0;
      10'h1ad: data = 32'h2c420030; // 004006b4: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h1ae: data = 32'h10400009; // 004006b8: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h1af: data = 32'h00000000; // 004006bc: SLL, REG[0]<=REG[0]<<0;
      10'h1b0: data = 32'h24020304; // 004006c0: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h1b1: data = 32'h8fc30008; // 004006c4: LW, REG[3]<=RAM[REG[30]+8];
      10'h1b2: data = 32'h00000000; // 004006c8: SLL, REG[0]<=REG[0]<<0;
      10'h1b3: data = 32'h8c630000; // 004006cc: LW, REG[3]<=RAM[REG[3]+0];
      10'h1b4: data = 32'h00000000; // 004006d0: SLL, REG[0]<=REG[0]<<0;
      10'h1b5: data = 32'hac430000; // 004006d4: SW, RAM[REG[2]+0]<=REG[3];
      10'h1b6: data = 32'h081001f1; // 004006d8: J, PC<=0x001001f1*4(=0x004007c4);
      10'h1b7: data = 32'h00000000; // 004006dc: SLL, REG[0]<=REG[0]<<0;
      10'h1b8: data = 32'h8fc20008; // 004006e0: LW, REG[2]<=RAM[REG[30]+8];
      10'h1b9: data = 32'h00000000; // 004006e4: SLL, REG[0]<=REG[0]<<0;
      10'h1ba: data = 32'h8c430000; // 004006e8: LW, REG[3]<=RAM[REG[2]+0];
      10'h1bb: data = 32'h2402003f; // 004006ec: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h1bc: data = 32'h14620006; // 004006f0: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1bd: data = 32'h00000000; // 004006f4: SLL, REG[0]<=REG[0]<<0;
      10'h1be: data = 32'h24030304; // 004006f8: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h1bf: data = 32'h2402003a; // 004006fc: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h1c0: data = 32'hac620000; // 00400700: SW, RAM[REG[3]+0]<=REG[2];
      10'h1c1: data = 32'h081001f1; // 00400704: J, PC<=0x001001f1*4(=0x004007c4);
      10'h1c2: data = 32'h00000000; // 00400708: SLL, REG[0]<=REG[0]<<0;
      10'h1c3: data = 32'h8fc20008; // 0040070c: LW, REG[2]<=RAM[REG[30]+8];
      10'h1c4: data = 32'h00000000; // 00400710: SLL, REG[0]<=REG[0]<<0;
      10'h1c5: data = 32'h8c430000; // 00400714: LW, REG[3]<=RAM[REG[2]+0];
      10'h1c6: data = 32'h2402003d; // 00400718: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h1c7: data = 32'h14620006; // 0040071c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1c8: data = 32'h00000000; // 00400720: SLL, REG[0]<=REG[0]<<0;
      10'h1c9: data = 32'h24030304; // 00400724: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h1ca: data = 32'h2402003b; // 00400728: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h1cb: data = 32'hac620000; // 0040072c: SW, RAM[REG[3]+0]<=REG[2];
      10'h1cc: data = 32'h081001f1; // 00400730: J, PC<=0x001001f1*4(=0x004007c4);
      10'h1cd: data = 32'h00000000; // 00400734: SLL, REG[0]<=REG[0]<<0;
      10'h1ce: data = 32'h8fc20008; // 00400738: LW, REG[2]<=RAM[REG[30]+8];
      10'h1cf: data = 32'h00000000; // 0040073c: SLL, REG[0]<=REG[0]<<0;
      10'h1d0: data = 32'h8c430000; // 00400740: LW, REG[3]<=RAM[REG[2]+0];
      10'h1d1: data = 32'h2402003b; // 00400744: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h1d2: data = 32'h14620006; // 00400748: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1d3: data = 32'h00000000; // 0040074c: SLL, REG[0]<=REG[0]<<0;
      10'h1d4: data = 32'h24030304; // 00400750: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h1d5: data = 32'h2402003c; // 00400754: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h1d6: data = 32'hac620000; // 00400758: SW, RAM[REG[3]+0]<=REG[2];
      10'h1d7: data = 32'h081001f1; // 0040075c: J, PC<=0x001001f1*4(=0x004007c4);
      10'h1d8: data = 32'h00000000; // 00400760: SLL, REG[0]<=REG[0]<<0;
      10'h1d9: data = 32'h8fc20008; // 00400764: LW, REG[2]<=RAM[REG[30]+8];
      10'h1da: data = 32'h00000000; // 00400768: SLL, REG[0]<=REG[0]<<0;
      10'h1db: data = 32'h8c430000; // 0040076c: LW, REG[3]<=RAM[REG[2]+0];
      10'h1dc: data = 32'h2402003a; // 00400770: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h1dd: data = 32'h14620006; // 00400774: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1de: data = 32'h00000000; // 00400778: SLL, REG[0]<=REG[0]<<0;
      10'h1df: data = 32'h24030304; // 0040077c: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h1e0: data = 32'h2402003d; // 00400780: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h1e1: data = 32'hac620000; // 00400784: SW, RAM[REG[3]+0]<=REG[2];
      10'h1e2: data = 32'h081001f1; // 00400788: J, PC<=0x001001f1*4(=0x004007c4);
      10'h1e3: data = 32'h00000000; // 0040078c: SLL, REG[0]<=REG[0]<<0;
      10'h1e4: data = 32'h8fc20008; // 00400790: LW, REG[2]<=RAM[REG[30]+8];
      10'h1e5: data = 32'h00000000; // 00400794: SLL, REG[0]<=REG[0]<<0;
      10'h1e6: data = 32'h8c430000; // 00400798: LW, REG[3]<=RAM[REG[2]+0];
      10'h1e7: data = 32'h2402000a; // 0040079c: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h1e8: data = 32'h14620006; // 004007a0: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1e9: data = 32'h00000000; // 004007a4: SLL, REG[0]<=REG[0]<<0;
      10'h1ea: data = 32'h24030304; // 004007a8: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h1eb: data = 32'h2402003e; // 004007ac: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h1ec: data = 32'hac620000; // 004007b0: SW, RAM[REG[3]+0]<=REG[2];
      10'h1ed: data = 32'h081001f1; // 004007b4: J, PC<=0x001001f1*4(=0x004007c4);
      10'h1ee: data = 32'h00000000; // 004007b8: SLL, REG[0]<=REG[0]<<0;
      10'h1ef: data = 32'h24020304; // 004007bc: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h1f0: data = 32'hac400000; // 004007c0: SW, RAM[REG[2]+0]<=REG[0];
      10'h1f1: data = 32'h24030300; // 004007c4: ADDIU, REG[3]<=REG[0]+768(=0x00000300);
      10'h1f2: data = 32'h24020001; // 004007c8: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h1f3: data = 32'hac620000; // 004007cc: SW, RAM[REG[3]+0]<=REG[2];
      10'h1f4: data = 32'h8fc20008; // 004007d0: LW, REG[2]<=RAM[REG[30]+8];
      10'h1f5: data = 32'h00000000; // 004007d4: SLL, REG[0]<=REG[0]<<0;
      10'h1f6: data = 32'h24420004; // 004007d8: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h1f7: data = 32'hafc20008; // 004007dc: SW, RAM[REG[30]+8]<=REG[2];
      10'h1f8: data = 32'h8fc20008; // 004007e0: LW, REG[2]<=RAM[REG[30]+8];
      10'h1f9: data = 32'h00000000; // 004007e4: SLL, REG[0]<=REG[0]<<0;
      10'h1fa: data = 32'h8c420000; // 004007e8: LW, REG[2]<=RAM[REG[2]+0];
      10'h1fb: data = 32'h00000000; // 004007ec: SLL, REG[0]<=REG[0]<<0;
      10'h1fc: data = 32'h1440ff3f; // 004007f0: BNE, PC<=(REG[2] != REG[0])?PC+4+65343*4:PC+4;
      10'h1fd: data = 32'h00000000; // 004007f4: SLL, REG[0]<=REG[0]<<0;
      10'h1fe: data = 32'h03c0e821; // 004007f8: ADDU, REG[29]<=REG[30]+REG[0];
      10'h1ff: data = 32'h8fbe0000; // 004007fc: LW, REG[30]<=RAM[REG[29]+0];
      10'h200: data = 32'h27bd0008; // 00400800: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h201: data = 32'h03e00008; // 00400804: JR, PC<=REG[31];
      10'h202: data = 32'h00000000; // 00400808: SLL, REG[0]<=REG[0]<<0;
      10'h203: data = 32'h00000000; // 0040080c: SLL, REG[0]<=REG[0]<<0;
    endcase
  end

  assign rom_data = data;
endmodule
